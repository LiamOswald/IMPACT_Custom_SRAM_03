VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO truncation_SRAM
  CLASS BLOCK ;
  FOREIGN truncation_SRAM ;
  ORIGIN 3.950 -17.900 ;
  SIZE 263.200 BY 2015.700 ;
  PIN DataOut31
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 241.400 17.900 241.700 19.900 ;
    END
  END DataOut31
  PIN DataOut30
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 240.100 17.900 240.400 19.900 ;
    END
  END DataOut30
  PIN DataOut29
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 238.800 17.900 239.100 19.900 ;
    END
  END DataOut29
  PIN DataOut28
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 237.500 17.900 237.800 19.900 ;
    END
  END DataOut28
  PIN DataOut27
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 215.100 17.900 215.400 19.900 ;
    END
  END DataOut27
  PIN DataOut26
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 213.800 17.900 214.100 19.900 ;
    END
  END DataOut26
  PIN DataOut25
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 212.500 17.900 212.800 19.900 ;
    END
  END DataOut25
  PIN DataOut24
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 211.200 17.900 211.500 19.900 ;
    END
  END DataOut24
  PIN DataOut23
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 181.000 17.900 181.300 19.900 ;
    END
  END DataOut23
  PIN DataOut22
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 179.700 17.900 180.000 19.900 ;
    END
  END DataOut22
  PIN DataOut21
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 178.400 17.900 178.700 19.900 ;
    END
  END DataOut21
  PIN DataOut20
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 177.100 17.900 177.400 19.900 ;
    END
  END DataOut20
  PIN DataOut19
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 154.700 17.900 155.000 19.900 ;
    END
  END DataOut19
  PIN DataOut18
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 153.400 17.900 153.700 19.900 ;
    END
  END DataOut18
  PIN DataOut17
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 152.100 17.900 152.400 19.900 ;
    END
  END DataOut17
  PIN DataOut16
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 150.800 17.900 151.100 19.900 ;
    END
  END DataOut16
  PIN DataOut15
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 120.600 17.900 120.900 19.900 ;
    END
  END DataOut15
  PIN DataOut14
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 119.300 17.900 119.600 19.900 ;
    END
  END DataOut14
  PIN DataOut13
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 118.000 17.900 118.300 19.900 ;
    END
  END DataOut13
  PIN DataOut12
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 116.700 17.900 117.000 19.900 ;
    END
  END DataOut12
  PIN DataOut11
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 94.300 17.900 94.600 19.900 ;
    END
  END DataOut11
  PIN DataOut10
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 93.000 17.900 93.300 19.900 ;
    END
  END DataOut10
  PIN DataOut9
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 91.700 17.900 92.000 19.900 ;
    END
  END DataOut9
  PIN DataOut8
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 90.400 17.900 90.700 19.900 ;
    END
  END DataOut8
  PIN DataOut7
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 60.200 17.900 60.500 19.900 ;
    END
  END DataOut7
  PIN DataOut6
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 58.900 17.900 59.200 19.900 ;
    END
  END DataOut6
  PIN DataOut5
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 57.600 17.900 57.900 19.900 ;
    END
  END DataOut5
  PIN DataOut4
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 56.300 17.900 56.600 19.900 ;
    END
  END DataOut4
  PIN DataOut3
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 33.900 17.900 34.200 19.900 ;
    END
  END DataOut3
  PIN DataOut2
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 32.600 17.900 32.900 19.900 ;
    END
  END DataOut2
  PIN DataOut1
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 31.300 17.900 31.600 19.900 ;
    END
  END DataOut1
  PIN DataOut0
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER met2 ;
        RECT 30.000 17.900 30.300 19.900 ;
    END
  END DataOut0
  PIN Trunk0
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 12.600 17.900 12.900 19.900 ;
    END
  END Trunk0
  PIN Trunk1
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 13.900 17.900 14.200 19.900 ;
    END
  END Trunk1
  PIN Trunk2
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 15.200 17.900 15.500 19.900 ;
    END
  END Trunk2
  PIN Trunk3
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 16.500 17.900 16.800 19.900 ;
    END
  END Trunk3
  PIN Trunk4
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 17.800 17.900 18.100 19.900 ;
    END
  END Trunk4
  PIN Trunk5
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 19.100 17.900 19.400 19.900 ;
    END
  END Trunk5
  PIN Trunk6
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 20.400 17.900 20.700 19.900 ;
    END
  END Trunk6
  PIN Trunk7
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 21.700 17.900 22.000 19.900 ;
    END
  END Trunk7
  PIN Trunk8
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 65.500 17.900 65.800 19.900 ;
    END
  END Trunk8
  PIN Trunk9
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 66.800 17.900 67.100 19.900 ;
    END
  END Trunk9
  PIN Trunk10
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 68.100 17.900 68.400 19.900 ;
    END
  END Trunk10
  PIN Trunk11
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 69.400 17.900 69.700 19.900 ;
    END
  END Trunk11
  PIN Trunk12
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 70.700 17.900 71.000 19.900 ;
    END
  END Trunk12
  PIN Trunk13
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 72.000 17.900 72.300 19.900 ;
    END
  END Trunk13
  PIN Trunk14
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 73.300 17.900 73.600 19.900 ;
    END
  END Trunk14
  PIN Trunk15
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 74.600 17.900 74.900 19.900 ;
    END
  END Trunk15
  PIN Trunk16
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 125.900 17.900 126.200 19.900 ;
    END
  END Trunk16
  PIN Trunk17
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 127.200 17.900 127.500 19.900 ;
    END
  END Trunk17
  PIN Trunk18
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 128.500 17.900 128.800 19.900 ;
    END
  END Trunk18
  PIN Trunk19
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 129.800 17.900 130.100 19.900 ;
    END
  END Trunk19
  PIN Trunk20
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 131.100 17.900 131.400 19.900 ;
    END
  END Trunk20
  PIN Trunk21
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 132.400 17.900 132.700 19.900 ;
    END
  END Trunk21
  PIN Trunk22
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 133.700 17.900 134.000 19.900 ;
    END
  END Trunk22
  PIN Trunk23
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 135.000 17.900 135.300 19.900 ;
    END
  END Trunk23
  PIN Trunk24
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 186.300 17.900 186.600 19.900 ;
    END
  END Trunk24
  PIN Trunk25
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 187.600 17.900 187.900 19.900 ;
    END
  END Trunk25
  PIN Trunk26
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 188.900 17.900 189.200 19.900 ;
    END
  END Trunk26
  PIN Trunk27
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 190.200 17.900 190.500 19.900 ;
    END
  END Trunk27
  PIN Trunk28
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 191.500 17.900 191.800 19.900 ;
    END
  END Trunk28
  PIN Trunk29
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 192.800 17.900 193.100 19.900 ;
    END
  END Trunk29
  PIN Trunk30
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 194.100 17.900 194.400 19.900 ;
    END
  END Trunk30
  PIN Trunk31
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 195.400 17.900 195.700 19.900 ;
    END
  END Trunk31
  PIN Tail_In
    ANTENNAGATEAREA 1.134000 ;
    PORT
      LAYER met2 ;
        RECT 233.400 17.900 233.700 19.900 ;
    END
  END Tail_In
  PIN vccd1
    ANTENNADIFFAREA 1498.728394 ;
    PORT
      LAYER met2 ;
        RECT -1.750 2031.600 0.250 2033.600 ;
        RECT 21.250 2031.600 21.800 2033.200 ;
        RECT 255.250 2031.600 257.250 2033.600 ;
      LAYER via2 ;
        RECT -1.250 2032.100 -0.250 2033.100 ;
        RECT 21.350 2032.000 21.700 2033.100 ;
        RECT 255.750 2032.100 256.750 2033.100 ;
      LAYER met3 ;
        RECT -3.950 2031.600 257.250 2033.600 ;
        RECT -3.950 19.900 257.250 21.900 ;
    END
  END vccd1
  PIN vssd1
    ANTENNADIFFAREA 8225.771484 ;
    PORT
      LAYER met3 ;
        RECT -3.950 2026.600 -1.950 2028.600 ;
        RECT -3.950 24.900 257.250 26.900 ;
    END
  END vssd1
  PIN Byte_Mode_EnableBar
    ANTENNAGATEAREA 1.512000 ;
    PORT
      LAYER met2 ;
        RECT 26.650 17.900 26.950 19.900 ;
    END
  END Byte_Mode_EnableBar
  PIN PRE
    ANTENNAGATEAREA 8.294400 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2021.850 -1.950 2022.050 ;
        RECT -3.750 2021.250 -1.750 2021.850 ;
        RECT -3.750 2021.050 -1.950 2021.250 ;
    END
  END PRE
  PIN writeen
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 149.950 -1.950 150.150 ;
        RECT -3.750 149.350 -1.750 149.950 ;
        RECT -3.750 149.150 -1.950 149.350 ;
    END
  END writeen
  PIN readen
    ANTENNAGATEAREA 7.257600 ;
    PORT
      LAYER met3 ;
        RECT -3.750 162.450 -1.950 162.650 ;
        RECT -3.750 161.850 -1.750 162.450 ;
        RECT -3.750 161.650 -1.950 161.850 ;
    END
  END readen
  PIN DataIn31
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 135.900 259.250 136.600 ;
    END
  END DataIn31
  PIN DataIn30
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 133.800 259.250 134.500 ;
    END
  END DataIn30
  PIN DataIn29
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 131.700 259.250 132.400 ;
    END
  END DataIn29
  PIN DataIn28
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 129.600 259.250 130.300 ;
    END
  END DataIn28
  PIN DataIn27
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 127.500 259.250 128.200 ;
    END
  END DataIn27
  PIN DataIn26
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 125.400 259.250 126.100 ;
    END
  END DataIn26
  PIN DataIn25
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 123.300 259.250 124.000 ;
    END
  END DataIn25
  PIN DataIn24
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 121.200 259.250 121.900 ;
    END
  END DataIn24
  PIN DataIn23
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 119.100 259.250 119.800 ;
    END
  END DataIn23
  PIN DataIn22
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 117.000 259.250 117.700 ;
    END
  END DataIn22
  PIN DataIn21
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 114.900 259.250 115.600 ;
    END
  END DataIn21
  PIN DataIn20
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 112.800 259.250 113.500 ;
    END
  END DataIn20
  PIN DataIn19
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 110.700 259.250 111.400 ;
    END
  END DataIn19
  PIN DataIn18
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 108.600 259.250 109.300 ;
    END
  END DataIn18
  PIN DataIn17
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 106.500 259.250 107.200 ;
    END
  END DataIn17
  PIN DataIn16
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 257.250 104.400 259.250 105.100 ;
    END
  END DataIn16
  PIN DataIn15
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 105.050 -1.950 105.100 ;
        RECT -3.750 104.450 -1.750 105.050 ;
        RECT -3.750 104.400 -1.950 104.450 ;
    END
  END DataIn15
  PIN DataIn14
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 107.150 -1.950 107.200 ;
        RECT -3.750 106.550 -1.750 107.150 ;
        RECT -3.750 106.500 -1.950 106.550 ;
    END
  END DataIn14
  PIN DataIn13
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 109.250 -1.950 109.300 ;
        RECT -3.750 108.650 -1.750 109.250 ;
        RECT -3.750 108.600 -1.950 108.650 ;
    END
  END DataIn13
  PIN DataIn12
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 111.350 -1.950 111.400 ;
        RECT -3.750 110.750 -1.750 111.350 ;
        RECT -3.750 110.700 -1.950 110.750 ;
    END
  END DataIn12
  PIN DataIn11
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 113.450 -1.950 113.500 ;
        RECT -3.750 112.850 -1.750 113.450 ;
        RECT -3.750 112.800 -1.950 112.850 ;
    END
  END DataIn11
  PIN DataIn10
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 115.550 -1.950 115.600 ;
        RECT -3.750 114.950 -1.750 115.550 ;
        RECT -3.750 114.900 -1.950 114.950 ;
    END
  END DataIn10
  PIN DataIn9
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 117.650 -1.950 117.700 ;
        RECT -3.750 117.050 -1.750 117.650 ;
        RECT -3.750 117.000 -1.950 117.050 ;
    END
  END DataIn9
  PIN DataIn8
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 119.750 -1.950 119.800 ;
        RECT -3.750 119.150 -1.750 119.750 ;
        RECT -3.750 119.100 -1.950 119.150 ;
    END
  END DataIn8
  PIN DataIn7
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 121.850 -1.950 121.900 ;
        RECT -3.750 121.250 -1.750 121.850 ;
        RECT -3.750 121.200 -1.950 121.250 ;
    END
  END DataIn7
  PIN DataIn6
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 123.950 -1.950 124.000 ;
        RECT -3.750 123.350 -1.750 123.950 ;
        RECT -3.750 123.300 -1.950 123.350 ;
    END
  END DataIn6
  PIN DataIn5
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 126.050 -1.950 126.100 ;
        RECT -3.750 125.450 -1.750 126.050 ;
        RECT -3.750 125.400 -1.950 125.450 ;
    END
  END DataIn5
  PIN DataIn4
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 128.150 -1.950 128.200 ;
        RECT -3.750 127.550 -1.750 128.150 ;
        RECT -3.750 127.500 -1.950 127.550 ;
    END
  END DataIn4
  PIN DataIn3
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 130.250 -1.950 130.300 ;
        RECT -3.750 129.650 -1.750 130.250 ;
        RECT -3.750 129.600 -1.950 129.650 ;
    END
  END DataIn3
  PIN DataIn2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 132.350 -1.950 132.400 ;
        RECT -3.750 131.750 -1.750 132.350 ;
        RECT -3.750 131.700 -1.950 131.750 ;
    END
  END DataIn2
  PIN DataIn1
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 134.450 -1.950 134.500 ;
        RECT -3.750 133.850 -1.750 134.450 ;
        RECT -3.750 133.800 -1.950 133.850 ;
    END
  END DataIn1
  PIN DataIn0
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 136.550 -1.950 136.600 ;
        RECT -3.750 135.950 -1.750 136.550 ;
        RECT -3.750 135.900 -1.950 135.950 ;
    END
  END DataIn0
  PIN WL0
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2016.650 -1.950 2016.850 ;
        RECT -3.750 2016.050 -1.750 2016.650 ;
        RECT -3.750 2015.850 -1.950 2016.050 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2015.300 -1.950 2015.500 ;
        RECT -3.750 2014.700 -1.750 2015.300 ;
        RECT -3.750 2014.500 -1.950 2014.700 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2013.050 -1.950 2013.250 ;
        RECT -3.750 2012.450 -1.750 2013.050 ;
        RECT -3.750 2012.250 -1.950 2012.450 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2011.700 -1.950 2011.900 ;
        RECT -3.750 2011.100 -1.750 2011.700 ;
        RECT -3.750 2010.900 -1.950 2011.100 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2009.450 -1.950 2009.650 ;
        RECT -3.750 2008.850 -1.750 2009.450 ;
        RECT -3.750 2008.650 -1.950 2008.850 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2008.100 -1.950 2008.300 ;
        RECT -3.750 2007.500 -1.750 2008.100 ;
        RECT -3.750 2007.300 -1.950 2007.500 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2005.850 -1.950 2006.050 ;
        RECT -3.750 2005.250 -1.750 2005.850 ;
        RECT -3.750 2005.050 -1.950 2005.250 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2004.500 -1.950 2004.700 ;
        RECT -3.750 2003.900 -1.750 2004.500 ;
        RECT -3.750 2003.700 -1.950 2003.900 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2002.250 -1.950 2002.450 ;
        RECT -3.750 2001.650 -1.750 2002.250 ;
        RECT -3.750 2001.450 -1.950 2001.650 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 2000.900 -1.950 2001.100 ;
        RECT -3.750 2000.300 -1.750 2000.900 ;
        RECT -3.750 2000.100 -1.950 2000.300 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1998.650 -1.950 1998.850 ;
        RECT -3.750 1998.050 -1.750 1998.650 ;
        RECT -3.750 1997.850 -1.950 1998.050 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1997.300 -1.950 1997.500 ;
        RECT -3.750 1996.700 -1.750 1997.300 ;
        RECT -3.750 1996.500 -1.950 1996.700 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1995.050 -1.950 1995.250 ;
        RECT -3.750 1994.450 -1.750 1995.050 ;
        RECT -3.750 1994.250 -1.950 1994.450 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1993.700 -1.950 1993.900 ;
        RECT -3.750 1993.100 -1.750 1993.700 ;
        RECT -3.750 1992.900 -1.950 1993.100 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1991.450 -1.950 1991.650 ;
        RECT -3.750 1990.850 -1.750 1991.450 ;
        RECT -3.750 1990.650 -1.950 1990.850 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1990.100 -1.950 1990.300 ;
        RECT -3.750 1989.500 -1.750 1990.100 ;
        RECT -3.750 1989.300 -1.950 1989.500 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1987.850 -1.950 1988.050 ;
        RECT -3.750 1987.250 -1.750 1987.850 ;
        RECT -3.750 1987.050 -1.950 1987.250 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1986.500 -1.950 1986.700 ;
        RECT -3.750 1985.900 -1.750 1986.500 ;
        RECT -3.750 1985.700 -1.950 1985.900 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1984.250 -1.950 1984.450 ;
        RECT -3.750 1983.650 -1.750 1984.250 ;
        RECT -3.750 1983.450 -1.950 1983.650 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1982.900 -1.950 1983.100 ;
        RECT -3.750 1982.300 -1.750 1982.900 ;
        RECT -3.750 1982.100 -1.950 1982.300 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1980.650 -1.950 1980.850 ;
        RECT -3.750 1980.050 -1.750 1980.650 ;
        RECT -3.750 1979.850 -1.950 1980.050 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1979.300 -1.950 1979.500 ;
        RECT -3.750 1978.700 -1.750 1979.300 ;
        RECT -3.750 1978.500 -1.950 1978.700 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1977.050 -1.950 1977.250 ;
        RECT -3.750 1976.450 -1.750 1977.050 ;
        RECT -3.750 1976.250 -1.950 1976.450 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1975.700 -1.950 1975.900 ;
        RECT -3.750 1975.100 -1.750 1975.700 ;
        RECT -3.750 1974.900 -1.950 1975.100 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1973.450 -1.950 1973.650 ;
        RECT -3.750 1972.850 -1.750 1973.450 ;
        RECT -3.750 1972.650 -1.950 1972.850 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1972.100 -1.950 1972.300 ;
        RECT -3.750 1971.500 -1.750 1972.100 ;
        RECT -3.750 1971.300 -1.950 1971.500 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1969.850 -1.950 1970.050 ;
        RECT -3.750 1969.250 -1.750 1969.850 ;
        RECT -3.750 1969.050 -1.950 1969.250 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1968.500 -1.950 1968.700 ;
        RECT -3.750 1967.900 -1.750 1968.500 ;
        RECT -3.750 1967.700 -1.950 1967.900 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1966.250 -1.950 1966.450 ;
        RECT -3.750 1965.650 -1.750 1966.250 ;
        RECT -3.750 1965.450 -1.950 1965.650 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1964.900 -1.950 1965.100 ;
        RECT -3.750 1964.300 -1.750 1964.900 ;
        RECT -3.750 1964.100 -1.950 1964.300 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1962.650 -1.950 1962.850 ;
        RECT -3.750 1962.050 -1.750 1962.650 ;
        RECT -3.750 1961.850 -1.950 1962.050 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1961.300 -1.950 1961.500 ;
        RECT -3.750 1960.700 -1.750 1961.300 ;
        RECT -3.750 1960.500 -1.950 1960.700 ;
    END
  END WL31
  PIN WL32
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1959.050 -1.950 1959.250 ;
        RECT -3.750 1958.450 -1.750 1959.050 ;
        RECT -3.750 1958.250 -1.950 1958.450 ;
    END
  END WL32
  PIN WL33
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1957.700 -1.950 1957.900 ;
        RECT -3.750 1957.100 -1.750 1957.700 ;
        RECT -3.750 1956.900 -1.950 1957.100 ;
    END
  END WL33
  PIN WL34
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1955.450 -1.950 1955.650 ;
        RECT -3.750 1954.850 -1.750 1955.450 ;
        RECT -3.750 1954.650 -1.950 1954.850 ;
    END
  END WL34
  PIN WL35
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1954.100 -1.950 1954.300 ;
        RECT -3.750 1953.500 -1.750 1954.100 ;
        RECT -3.750 1953.300 -1.950 1953.500 ;
    END
  END WL35
  PIN WL36
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1951.850 -1.950 1952.050 ;
        RECT -3.750 1951.250 -1.750 1951.850 ;
        RECT -3.750 1951.050 -1.950 1951.250 ;
    END
  END WL36
  PIN WL37
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1950.500 -1.950 1950.700 ;
        RECT -3.750 1949.900 -1.750 1950.500 ;
        RECT -3.750 1949.700 -1.950 1949.900 ;
    END
  END WL37
  PIN WL38
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1948.250 -1.950 1948.450 ;
        RECT -3.750 1947.650 -1.750 1948.250 ;
        RECT -3.750 1947.450 -1.950 1947.650 ;
    END
  END WL38
  PIN WL39
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1946.900 -1.950 1947.100 ;
        RECT -3.750 1946.300 -1.750 1946.900 ;
        RECT -3.750 1946.100 -1.950 1946.300 ;
    END
  END WL39
  PIN WL40
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1944.650 -1.950 1944.850 ;
        RECT -3.750 1944.050 -1.750 1944.650 ;
        RECT -3.750 1943.850 -1.950 1944.050 ;
    END
  END WL40
  PIN WL41
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1943.300 -1.950 1943.500 ;
        RECT -3.750 1942.700 -1.750 1943.300 ;
        RECT -3.750 1942.500 -1.950 1942.700 ;
    END
  END WL41
  PIN WL42
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1941.050 -1.950 1941.250 ;
        RECT -3.750 1940.450 -1.750 1941.050 ;
        RECT -3.750 1940.250 -1.950 1940.450 ;
    END
  END WL42
  PIN WL43
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1939.700 -1.950 1939.900 ;
        RECT -3.750 1939.100 -1.750 1939.700 ;
        RECT -3.750 1938.900 -1.950 1939.100 ;
    END
  END WL43
  PIN WL44
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1937.450 -1.950 1937.650 ;
        RECT -3.750 1936.850 -1.750 1937.450 ;
        RECT -3.750 1936.650 -1.950 1936.850 ;
    END
  END WL44
  PIN WL45
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1936.100 -1.950 1936.300 ;
        RECT -3.750 1935.500 -1.750 1936.100 ;
        RECT -3.750 1935.300 -1.950 1935.500 ;
    END
  END WL45
  PIN WL46
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1933.850 -1.950 1934.050 ;
        RECT -3.750 1933.250 -1.750 1933.850 ;
        RECT -3.750 1933.050 -1.950 1933.250 ;
    END
  END WL46
  PIN WL47
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1932.500 -1.950 1932.700 ;
        RECT -3.750 1931.900 -1.750 1932.500 ;
        RECT -3.750 1931.700 -1.950 1931.900 ;
    END
  END WL47
  PIN WL48
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1930.250 -1.950 1930.450 ;
        RECT -3.750 1929.650 -1.750 1930.250 ;
        RECT -3.750 1929.450 -1.950 1929.650 ;
    END
  END WL48
  PIN WL49
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1928.900 -1.950 1929.100 ;
        RECT -3.750 1928.300 -1.750 1928.900 ;
        RECT -3.750 1928.100 -1.950 1928.300 ;
    END
  END WL49
  PIN WL50
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1926.650 -1.950 1926.850 ;
        RECT -3.750 1926.050 -1.750 1926.650 ;
        RECT -3.750 1925.850 -1.950 1926.050 ;
    END
  END WL50
  PIN WL51
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1925.300 -1.950 1925.500 ;
        RECT -3.750 1924.700 -1.750 1925.300 ;
        RECT -3.750 1924.500 -1.950 1924.700 ;
    END
  END WL51
  PIN WL52
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1923.050 -1.950 1923.250 ;
        RECT -3.750 1922.450 -1.750 1923.050 ;
        RECT -3.750 1922.250 -1.950 1922.450 ;
    END
  END WL52
  PIN WL53
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1921.700 -1.950 1921.900 ;
        RECT -3.750 1921.100 -1.750 1921.700 ;
        RECT -3.750 1920.900 -1.950 1921.100 ;
    END
  END WL53
  PIN WL54
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1919.450 -1.950 1919.650 ;
        RECT -3.750 1918.850 -1.750 1919.450 ;
        RECT -3.750 1918.650 -1.950 1918.850 ;
    END
  END WL54
  PIN WL55
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1918.100 -1.950 1918.300 ;
        RECT -3.750 1917.500 -1.750 1918.100 ;
        RECT -3.750 1917.300 -1.950 1917.500 ;
    END
  END WL55
  PIN WL56
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1915.850 -1.950 1916.050 ;
        RECT -3.750 1915.250 -1.750 1915.850 ;
        RECT -3.750 1915.050 -1.950 1915.250 ;
    END
  END WL56
  PIN WL57
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1914.500 -1.950 1914.700 ;
        RECT -3.750 1913.900 -1.750 1914.500 ;
        RECT -3.750 1913.700 -1.950 1913.900 ;
    END
  END WL57
  PIN WL58
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1912.250 -1.950 1912.450 ;
        RECT -3.750 1911.650 -1.750 1912.250 ;
        RECT -3.750 1911.450 -1.950 1911.650 ;
    END
  END WL58
  PIN WL59
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1910.900 -1.950 1911.100 ;
        RECT -3.750 1910.300 -1.750 1910.900 ;
        RECT -3.750 1910.100 -1.950 1910.300 ;
    END
  END WL59
  PIN WL60
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1908.650 -1.950 1908.850 ;
        RECT -3.750 1908.050 -1.750 1908.650 ;
        RECT -3.750 1907.850 -1.950 1908.050 ;
    END
  END WL60
  PIN WL61
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1907.300 -1.950 1907.500 ;
        RECT -3.750 1906.700 -1.750 1907.300 ;
        RECT -3.750 1906.500 -1.950 1906.700 ;
    END
  END WL61
  PIN WL62
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1905.050 -1.950 1905.250 ;
        RECT -3.750 1904.450 -1.750 1905.050 ;
        RECT -3.750 1904.250 -1.950 1904.450 ;
    END
  END WL62
  PIN WL63
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1903.700 -1.950 1903.900 ;
        RECT -3.750 1903.100 -1.750 1903.700 ;
        RECT -3.750 1902.900 -1.950 1903.100 ;
    END
  END WL63
  PIN WL64
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1901.450 -1.950 1901.650 ;
        RECT -3.750 1900.850 -1.750 1901.450 ;
        RECT -3.750 1900.650 -1.950 1900.850 ;
    END
  END WL64
  PIN WL65
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1900.100 -1.950 1900.300 ;
        RECT -3.750 1899.500 -1.750 1900.100 ;
        RECT -3.750 1899.300 -1.950 1899.500 ;
    END
  END WL65
  PIN WL66
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1897.850 -1.950 1898.050 ;
        RECT -3.750 1897.250 -1.750 1897.850 ;
        RECT -3.750 1897.050 -1.950 1897.250 ;
    END
  END WL66
  PIN WL67
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1896.500 -1.950 1896.700 ;
        RECT -3.750 1895.900 -1.750 1896.500 ;
        RECT -3.750 1895.700 -1.950 1895.900 ;
    END
  END WL67
  PIN WL68
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1894.250 -1.950 1894.450 ;
        RECT -3.750 1893.650 -1.750 1894.250 ;
        RECT -3.750 1893.450 -1.950 1893.650 ;
    END
  END WL68
  PIN WL69
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1892.900 -1.950 1893.100 ;
        RECT -3.750 1892.300 -1.750 1892.900 ;
        RECT -3.750 1892.100 -1.950 1892.300 ;
    END
  END WL69
  PIN WL70
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1890.650 -1.950 1890.850 ;
        RECT -3.750 1890.050 -1.750 1890.650 ;
        RECT -3.750 1889.850 -1.950 1890.050 ;
    END
  END WL70
  PIN WL71
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1889.300 -1.950 1889.500 ;
        RECT -3.750 1888.700 -1.750 1889.300 ;
        RECT -3.750 1888.500 -1.950 1888.700 ;
    END
  END WL71
  PIN WL72
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1887.050 -1.950 1887.250 ;
        RECT -3.750 1886.450 -1.750 1887.050 ;
        RECT -3.750 1886.250 -1.950 1886.450 ;
    END
  END WL72
  PIN WL73
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1885.700 -1.950 1885.900 ;
        RECT -3.750 1885.100 -1.750 1885.700 ;
        RECT -3.750 1884.900 -1.950 1885.100 ;
    END
  END WL73
  PIN WL74
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1883.450 -1.950 1883.650 ;
        RECT -3.750 1882.850 -1.750 1883.450 ;
        RECT -3.750 1882.650 -1.950 1882.850 ;
    END
  END WL74
  PIN WL75
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1882.100 -1.950 1882.300 ;
        RECT -3.750 1881.500 -1.750 1882.100 ;
        RECT -3.750 1881.300 -1.950 1881.500 ;
    END
  END WL75
  PIN WL76
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1879.850 -1.950 1880.050 ;
        RECT -3.750 1879.250 -1.750 1879.850 ;
        RECT -3.750 1879.050 -1.950 1879.250 ;
    END
  END WL76
  PIN WL77
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1878.500 -1.950 1878.700 ;
        RECT -3.750 1877.900 -1.750 1878.500 ;
        RECT -3.750 1877.700 -1.950 1877.900 ;
    END
  END WL77
  PIN WL78
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1876.250 -1.950 1876.450 ;
        RECT -3.750 1875.650 -1.750 1876.250 ;
        RECT -3.750 1875.450 -1.950 1875.650 ;
    END
  END WL78
  PIN WL79
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1874.900 -1.950 1875.100 ;
        RECT -3.750 1874.300 -1.750 1874.900 ;
        RECT -3.750 1874.100 -1.950 1874.300 ;
    END
  END WL79
  PIN WL80
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1872.650 -1.950 1872.850 ;
        RECT -3.750 1872.050 -1.750 1872.650 ;
        RECT -3.750 1871.850 -1.950 1872.050 ;
    END
  END WL80
  PIN WL81
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1871.300 -1.950 1871.500 ;
        RECT -3.750 1870.700 -1.750 1871.300 ;
        RECT -3.750 1870.500 -1.950 1870.700 ;
    END
  END WL81
  PIN WL82
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1869.050 -1.950 1869.250 ;
        RECT -3.750 1868.450 -1.750 1869.050 ;
        RECT -3.750 1868.250 -1.950 1868.450 ;
    END
  END WL82
  PIN WL83
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1867.700 -1.950 1867.900 ;
        RECT -3.750 1867.100 -1.750 1867.700 ;
        RECT -3.750 1866.900 -1.950 1867.100 ;
    END
  END WL83
  PIN WL84
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1865.450 -1.950 1865.650 ;
        RECT -3.750 1864.850 -1.750 1865.450 ;
        RECT -3.750 1864.650 -1.950 1864.850 ;
    END
  END WL84
  PIN WL85
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1864.100 -1.950 1864.300 ;
        RECT -3.750 1863.500 -1.750 1864.100 ;
        RECT -3.750 1863.300 -1.950 1863.500 ;
    END
  END WL85
  PIN WL86
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1861.850 -1.950 1862.050 ;
        RECT -3.750 1861.250 -1.750 1861.850 ;
        RECT -3.750 1861.050 -1.950 1861.250 ;
    END
  END WL86
  PIN WL87
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1860.500 -1.950 1860.700 ;
        RECT -3.750 1859.900 -1.750 1860.500 ;
        RECT -3.750 1859.700 -1.950 1859.900 ;
    END
  END WL87
  PIN WL88
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1858.250 -1.950 1858.450 ;
        RECT -3.750 1857.650 -1.750 1858.250 ;
        RECT -3.750 1857.450 -1.950 1857.650 ;
    END
  END WL88
  PIN WL89
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1856.900 -1.950 1857.100 ;
        RECT -3.750 1856.300 -1.750 1856.900 ;
        RECT -3.750 1856.100 -1.950 1856.300 ;
    END
  END WL89
  PIN WL90
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1854.650 -1.950 1854.850 ;
        RECT -3.750 1854.050 -1.750 1854.650 ;
        RECT -3.750 1853.850 -1.950 1854.050 ;
    END
  END WL90
  PIN WL91
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1853.300 -1.950 1853.500 ;
        RECT -3.750 1852.700 -1.750 1853.300 ;
        RECT -3.750 1852.500 -1.950 1852.700 ;
    END
  END WL91
  PIN WL92
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1851.050 -1.950 1851.250 ;
        RECT -3.750 1850.450 -1.750 1851.050 ;
        RECT -3.750 1850.250 -1.950 1850.450 ;
    END
  END WL92
  PIN WL93
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1849.700 -1.950 1849.900 ;
        RECT -3.750 1849.100 -1.750 1849.700 ;
        RECT -3.750 1848.900 -1.950 1849.100 ;
    END
  END WL93
  PIN WL94
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1847.450 -1.950 1847.650 ;
        RECT -3.750 1846.850 -1.750 1847.450 ;
        RECT -3.750 1846.650 -1.950 1846.850 ;
    END
  END WL94
  PIN WL95
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1846.100 -1.950 1846.300 ;
        RECT -3.750 1845.500 -1.750 1846.100 ;
        RECT -3.750 1845.300 -1.950 1845.500 ;
    END
  END WL95
  PIN WL96
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1843.850 -1.950 1844.050 ;
        RECT -3.750 1843.250 -1.750 1843.850 ;
        RECT -3.750 1843.050 -1.950 1843.250 ;
    END
  END WL96
  PIN WL97
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1842.500 -1.950 1842.700 ;
        RECT -3.750 1841.900 -1.750 1842.500 ;
        RECT -3.750 1841.700 -1.950 1841.900 ;
    END
  END WL97
  PIN WL98
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1840.250 -1.950 1840.450 ;
        RECT -3.750 1839.650 -1.750 1840.250 ;
        RECT -3.750 1839.450 -1.950 1839.650 ;
    END
  END WL98
  PIN WL99
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1838.900 -1.950 1839.100 ;
        RECT -3.750 1838.300 -1.750 1838.900 ;
        RECT -3.750 1838.100 -1.950 1838.300 ;
    END
  END WL99
  PIN WL100
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1836.650 -1.950 1836.850 ;
        RECT -3.750 1836.050 -1.750 1836.650 ;
        RECT -3.750 1835.850 -1.950 1836.050 ;
    END
  END WL100
  PIN WL101
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1835.300 -1.950 1835.500 ;
        RECT -3.750 1834.700 -1.750 1835.300 ;
        RECT -3.750 1834.500 -1.950 1834.700 ;
    END
  END WL101
  PIN WL102
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1833.050 -1.950 1833.250 ;
        RECT -3.750 1832.450 -1.750 1833.050 ;
        RECT -3.750 1832.250 -1.950 1832.450 ;
    END
  END WL102
  PIN WL103
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1831.700 -1.950 1831.900 ;
        RECT -3.750 1831.100 -1.750 1831.700 ;
        RECT -3.750 1830.900 -1.950 1831.100 ;
    END
  END WL103
  PIN WL104
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1829.450 -1.950 1829.650 ;
        RECT -3.750 1828.850 -1.750 1829.450 ;
        RECT -3.750 1828.650 -1.950 1828.850 ;
    END
  END WL104
  PIN WL105
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1828.100 -1.950 1828.300 ;
        RECT -3.750 1827.500 -1.750 1828.100 ;
        RECT -3.750 1827.300 -1.950 1827.500 ;
    END
  END WL105
  PIN WL106
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1825.850 -1.950 1826.050 ;
        RECT -3.750 1825.250 -1.750 1825.850 ;
        RECT -3.750 1825.050 -1.950 1825.250 ;
    END
  END WL106
  PIN WL107
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1824.500 -1.950 1824.700 ;
        RECT -3.750 1823.900 -1.750 1824.500 ;
        RECT -3.750 1823.700 -1.950 1823.900 ;
    END
  END WL107
  PIN WL108
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1822.250 -1.950 1822.450 ;
        RECT -3.750 1821.650 -1.750 1822.250 ;
        RECT -3.750 1821.450 -1.950 1821.650 ;
    END
  END WL108
  PIN WL109
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1820.900 -1.950 1821.100 ;
        RECT -3.750 1820.300 -1.750 1820.900 ;
        RECT -3.750 1820.100 -1.950 1820.300 ;
    END
  END WL109
  PIN WL110
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1818.650 -1.950 1818.850 ;
        RECT -3.750 1818.050 -1.750 1818.650 ;
        RECT -3.750 1817.850 -1.950 1818.050 ;
    END
  END WL110
  PIN WL111
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1817.300 -1.950 1817.500 ;
        RECT -3.750 1816.700 -1.750 1817.300 ;
        RECT -3.750 1816.500 -1.950 1816.700 ;
    END
  END WL111
  PIN WL112
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1815.050 -1.950 1815.250 ;
        RECT -3.750 1814.450 -1.750 1815.050 ;
        RECT -3.750 1814.250 -1.950 1814.450 ;
    END
  END WL112
  PIN WL113
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1813.700 -1.950 1813.900 ;
        RECT -3.750 1813.100 -1.750 1813.700 ;
        RECT -3.750 1812.900 -1.950 1813.100 ;
    END
  END WL113
  PIN WL114
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1810.900 -1.950 1811.100 ;
        RECT -3.750 1810.300 -1.750 1810.900 ;
        RECT -3.750 1810.100 -1.950 1810.300 ;
    END
  END WL114
  PIN WL115
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1809.550 -1.950 1809.750 ;
        RECT -3.750 1808.950 -1.750 1809.550 ;
        RECT -3.750 1808.750 -1.950 1808.950 ;
    END
  END WL115
  PIN WL116
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1807.300 -1.950 1807.500 ;
        RECT -3.750 1806.700 -1.750 1807.300 ;
        RECT -3.750 1806.500 -1.950 1806.700 ;
    END
  END WL116
  PIN WL117
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1805.950 -1.950 1806.150 ;
        RECT -3.750 1805.350 -1.750 1805.950 ;
        RECT -3.750 1805.150 -1.950 1805.350 ;
    END
  END WL117
  PIN WL118
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1803.700 -1.950 1803.900 ;
        RECT -3.750 1803.100 -1.750 1803.700 ;
        RECT -3.750 1802.900 -1.950 1803.100 ;
    END
  END WL118
  PIN WL119
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1802.350 -1.950 1802.550 ;
        RECT -3.750 1801.750 -1.750 1802.350 ;
        RECT -3.750 1801.550 -1.950 1801.750 ;
    END
  END WL119
  PIN WL120
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1800.100 -1.950 1800.300 ;
        RECT -3.750 1799.500 -1.750 1800.100 ;
        RECT -3.750 1799.300 -1.950 1799.500 ;
    END
  END WL120
  PIN WL121
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1798.750 -1.950 1798.950 ;
        RECT -3.750 1798.150 -1.750 1798.750 ;
        RECT -3.750 1797.950 -1.950 1798.150 ;
    END
  END WL121
  PIN WL122
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1796.500 -1.950 1796.700 ;
        RECT -3.750 1795.900 -1.750 1796.500 ;
        RECT -3.750 1795.700 -1.950 1795.900 ;
    END
  END WL122
  PIN WL123
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1795.150 -1.950 1795.350 ;
        RECT -3.750 1794.550 -1.750 1795.150 ;
        RECT -3.750 1794.350 -1.950 1794.550 ;
    END
  END WL123
  PIN WL124
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1792.900 -1.950 1793.100 ;
        RECT -3.750 1792.300 -1.750 1792.900 ;
        RECT -3.750 1792.100 -1.950 1792.300 ;
    END
  END WL124
  PIN WL125
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1791.550 -1.950 1791.750 ;
        RECT -3.750 1790.950 -1.750 1791.550 ;
        RECT -3.750 1790.750 -1.950 1790.950 ;
    END
  END WL125
  PIN WL126
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1789.300 -1.950 1789.500 ;
        RECT -3.750 1788.700 -1.750 1789.300 ;
        RECT -3.750 1788.500 -1.950 1788.700 ;
    END
  END WL126
  PIN WL127
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1787.950 -1.950 1788.150 ;
        RECT -3.750 1787.350 -1.750 1787.950 ;
        RECT -3.750 1787.150 -1.950 1787.350 ;
    END
  END WL127
  PIN WL128
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1785.700 -1.950 1785.900 ;
        RECT -3.750 1785.100 -1.750 1785.700 ;
        RECT -3.750 1784.900 -1.950 1785.100 ;
    END
  END WL128
  PIN WL129
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1784.350 -1.950 1784.550 ;
        RECT -3.750 1783.750 -1.750 1784.350 ;
        RECT -3.750 1783.550 -1.950 1783.750 ;
    END
  END WL129
  PIN WL130
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1782.100 -1.950 1782.300 ;
        RECT -3.750 1781.500 -1.750 1782.100 ;
        RECT -3.750 1781.300 -1.950 1781.500 ;
    END
  END WL130
  PIN WL131
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1780.750 -1.950 1780.950 ;
        RECT -3.750 1780.150 -1.750 1780.750 ;
        RECT -3.750 1779.950 -1.950 1780.150 ;
    END
  END WL131
  PIN WL132
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1778.500 -1.950 1778.700 ;
        RECT -3.750 1777.900 -1.750 1778.500 ;
        RECT -3.750 1777.700 -1.950 1777.900 ;
    END
  END WL132
  PIN WL133
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1777.150 -1.950 1777.350 ;
        RECT -3.750 1776.550 -1.750 1777.150 ;
        RECT -3.750 1776.350 -1.950 1776.550 ;
    END
  END WL133
  PIN WL134
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1774.900 -1.950 1775.100 ;
        RECT -3.750 1774.300 -1.750 1774.900 ;
        RECT -3.750 1774.100 -1.950 1774.300 ;
    END
  END WL134
  PIN WL135
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1773.550 -1.950 1773.750 ;
        RECT -3.750 1772.950 -1.750 1773.550 ;
        RECT -3.750 1772.750 -1.950 1772.950 ;
    END
  END WL135
  PIN WL136
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1771.300 -1.950 1771.500 ;
        RECT -3.750 1770.700 -1.750 1771.300 ;
        RECT -3.750 1770.500 -1.950 1770.700 ;
    END
  END WL136
  PIN WL137
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1769.950 -1.950 1770.150 ;
        RECT -3.750 1769.350 -1.750 1769.950 ;
        RECT -3.750 1769.150 -1.950 1769.350 ;
    END
  END WL137
  PIN WL138
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1767.700 -1.950 1767.900 ;
        RECT -3.750 1767.100 -1.750 1767.700 ;
        RECT -3.750 1766.900 -1.950 1767.100 ;
    END
  END WL138
  PIN WL139
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1766.350 -1.950 1766.550 ;
        RECT -3.750 1765.750 -1.750 1766.350 ;
        RECT -3.750 1765.550 -1.950 1765.750 ;
    END
  END WL139
  PIN WL140
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1764.100 -1.950 1764.300 ;
        RECT -3.750 1763.500 -1.750 1764.100 ;
        RECT -3.750 1763.300 -1.950 1763.500 ;
    END
  END WL140
  PIN WL141
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1762.750 -1.950 1762.950 ;
        RECT -3.750 1762.150 -1.750 1762.750 ;
        RECT -3.750 1761.950 -1.950 1762.150 ;
    END
  END WL141
  PIN WL142
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1760.500 -1.950 1760.700 ;
        RECT -3.750 1759.900 -1.750 1760.500 ;
        RECT -3.750 1759.700 -1.950 1759.900 ;
    END
  END WL142
  PIN WL143
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1759.150 -1.950 1759.350 ;
        RECT -3.750 1758.550 -1.750 1759.150 ;
        RECT -3.750 1758.350 -1.950 1758.550 ;
    END
  END WL143
  PIN WL144
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1756.900 -1.950 1757.100 ;
        RECT -3.750 1756.300 -1.750 1756.900 ;
        RECT -3.750 1756.100 -1.950 1756.300 ;
    END
  END WL144
  PIN WL145
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1755.550 -1.950 1755.750 ;
        RECT -3.750 1754.950 -1.750 1755.550 ;
        RECT -3.750 1754.750 -1.950 1754.950 ;
    END
  END WL145
  PIN WL146
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1753.300 -1.950 1753.500 ;
        RECT -3.750 1752.700 -1.750 1753.300 ;
        RECT -3.750 1752.500 -1.950 1752.700 ;
    END
  END WL146
  PIN WL147
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1751.950 -1.950 1752.150 ;
        RECT -3.750 1751.350 -1.750 1751.950 ;
        RECT -3.750 1751.150 -1.950 1751.350 ;
    END
  END WL147
  PIN WL148
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1749.700 -1.950 1749.900 ;
        RECT -3.750 1749.100 -1.750 1749.700 ;
        RECT -3.750 1748.900 -1.950 1749.100 ;
    END
  END WL148
  PIN WL149
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1748.350 -1.950 1748.550 ;
        RECT -3.750 1747.750 -1.750 1748.350 ;
        RECT -3.750 1747.550 -1.950 1747.750 ;
    END
  END WL149
  PIN WL150
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1746.100 -1.950 1746.300 ;
        RECT -3.750 1745.500 -1.750 1746.100 ;
        RECT -3.750 1745.300 -1.950 1745.500 ;
    END
  END WL150
  PIN WL151
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1744.750 -1.950 1744.950 ;
        RECT -3.750 1744.150 -1.750 1744.750 ;
        RECT -3.750 1743.950 -1.950 1744.150 ;
    END
  END WL151
  PIN WL152
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1742.500 -1.950 1742.700 ;
        RECT -3.750 1741.900 -1.750 1742.500 ;
        RECT -3.750 1741.700 -1.950 1741.900 ;
    END
  END WL152
  PIN WL153
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1741.150 -1.950 1741.350 ;
        RECT -3.750 1740.550 -1.750 1741.150 ;
        RECT -3.750 1740.350 -1.950 1740.550 ;
    END
  END WL153
  PIN WL154
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1738.900 -1.950 1739.100 ;
        RECT -3.750 1738.300 -1.750 1738.900 ;
        RECT -3.750 1738.100 -1.950 1738.300 ;
    END
  END WL154
  PIN WL155
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1737.550 -1.950 1737.750 ;
        RECT -3.750 1736.950 -1.750 1737.550 ;
        RECT -3.750 1736.750 -1.950 1736.950 ;
    END
  END WL155
  PIN WL156
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1735.300 -1.950 1735.500 ;
        RECT -3.750 1734.700 -1.750 1735.300 ;
        RECT -3.750 1734.500 -1.950 1734.700 ;
    END
  END WL156
  PIN WL157
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1733.950 -1.950 1734.150 ;
        RECT -3.750 1733.350 -1.750 1733.950 ;
        RECT -3.750 1733.150 -1.950 1733.350 ;
    END
  END WL157
  PIN WL158
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1731.700 -1.950 1731.900 ;
        RECT -3.750 1731.100 -1.750 1731.700 ;
        RECT -3.750 1730.900 -1.950 1731.100 ;
    END
  END WL158
  PIN WL159
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1730.350 -1.950 1730.550 ;
        RECT -3.750 1729.750 -1.750 1730.350 ;
        RECT -3.750 1729.550 -1.950 1729.750 ;
    END
  END WL159
  PIN WL160
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1728.100 -1.950 1728.300 ;
        RECT -3.750 1727.500 -1.750 1728.100 ;
        RECT -3.750 1727.300 -1.950 1727.500 ;
    END
  END WL160
  PIN WL161
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1726.750 -1.950 1726.950 ;
        RECT -3.750 1726.150 -1.750 1726.750 ;
        RECT -3.750 1725.950 -1.950 1726.150 ;
    END
  END WL161
  PIN WL162
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1724.500 -1.950 1724.700 ;
        RECT -3.750 1723.900 -1.750 1724.500 ;
        RECT -3.750 1723.700 -1.950 1723.900 ;
    END
  END WL162
  PIN WL163
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1723.150 -1.950 1723.350 ;
        RECT -3.750 1722.550 -1.750 1723.150 ;
        RECT -3.750 1722.350 -1.950 1722.550 ;
    END
  END WL163
  PIN WL164
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1720.900 -1.950 1721.100 ;
        RECT -3.750 1720.300 -1.750 1720.900 ;
        RECT -3.750 1720.100 -1.950 1720.300 ;
    END
  END WL164
  PIN WL165
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1719.550 -1.950 1719.750 ;
        RECT -3.750 1718.950 -1.750 1719.550 ;
        RECT -3.750 1718.750 -1.950 1718.950 ;
    END
  END WL165
  PIN WL166
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1717.300 -1.950 1717.500 ;
        RECT -3.750 1716.700 -1.750 1717.300 ;
        RECT -3.750 1716.500 -1.950 1716.700 ;
    END
  END WL166
  PIN WL167
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1715.950 -1.950 1716.150 ;
        RECT -3.750 1715.350 -1.750 1715.950 ;
        RECT -3.750 1715.150 -1.950 1715.350 ;
    END
  END WL167
  PIN WL168
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1713.700 -1.950 1713.900 ;
        RECT -3.750 1713.100 -1.750 1713.700 ;
        RECT -3.750 1712.900 -1.950 1713.100 ;
    END
  END WL168
  PIN WL169
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1712.350 -1.950 1712.550 ;
        RECT -3.750 1711.750 -1.750 1712.350 ;
        RECT -3.750 1711.550 -1.950 1711.750 ;
    END
  END WL169
  PIN WL170
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1710.100 -1.950 1710.300 ;
        RECT -3.750 1709.500 -1.750 1710.100 ;
        RECT -3.750 1709.300 -1.950 1709.500 ;
    END
  END WL170
  PIN WL171
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1708.750 -1.950 1708.950 ;
        RECT -3.750 1708.150 -1.750 1708.750 ;
        RECT -3.750 1707.950 -1.950 1708.150 ;
    END
  END WL171
  PIN WL172
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1706.500 -1.950 1706.700 ;
        RECT -3.750 1705.900 -1.750 1706.500 ;
        RECT -3.750 1705.700 -1.950 1705.900 ;
    END
  END WL172
  PIN WL173
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1705.150 -1.950 1705.350 ;
        RECT -3.750 1704.550 -1.750 1705.150 ;
        RECT -3.750 1704.350 -1.950 1704.550 ;
    END
  END WL173
  PIN WL174
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1702.900 -1.950 1703.100 ;
        RECT -3.750 1702.300 -1.750 1702.900 ;
        RECT -3.750 1702.100 -1.950 1702.300 ;
    END
  END WL174
  PIN WL175
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1701.550 -1.950 1701.750 ;
        RECT -3.750 1700.950 -1.750 1701.550 ;
        RECT -3.750 1700.750 -1.950 1700.950 ;
    END
  END WL175
  PIN WL176
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1699.300 -1.950 1699.500 ;
        RECT -3.750 1698.700 -1.750 1699.300 ;
        RECT -3.750 1698.500 -1.950 1698.700 ;
    END
  END WL176
  PIN WL177
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1697.950 -1.950 1698.150 ;
        RECT -3.750 1697.350 -1.750 1697.950 ;
        RECT -3.750 1697.150 -1.950 1697.350 ;
    END
  END WL177
  PIN WL178
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1695.700 -1.950 1695.900 ;
        RECT -3.750 1695.100 -1.750 1695.700 ;
        RECT -3.750 1694.900 -1.950 1695.100 ;
    END
  END WL178
  PIN WL179
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1694.350 -1.950 1694.550 ;
        RECT -3.750 1693.750 -1.750 1694.350 ;
        RECT -3.750 1693.550 -1.950 1693.750 ;
    END
  END WL179
  PIN WL180
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1692.100 -1.950 1692.300 ;
        RECT -3.750 1691.500 -1.750 1692.100 ;
        RECT -3.750 1691.300 -1.950 1691.500 ;
    END
  END WL180
  PIN WL181
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1690.750 -1.950 1690.950 ;
        RECT -3.750 1690.150 -1.750 1690.750 ;
        RECT -3.750 1689.950 -1.950 1690.150 ;
    END
  END WL181
  PIN WL182
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1688.500 -1.950 1688.700 ;
        RECT -3.750 1687.900 -1.750 1688.500 ;
        RECT -3.750 1687.700 -1.950 1687.900 ;
    END
  END WL182
  PIN WL183
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1687.150 -1.950 1687.350 ;
        RECT -3.750 1686.550 -1.750 1687.150 ;
        RECT -3.750 1686.350 -1.950 1686.550 ;
    END
  END WL183
  PIN WL184
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1684.900 -1.950 1685.100 ;
        RECT -3.750 1684.300 -1.750 1684.900 ;
        RECT -3.750 1684.100 -1.950 1684.300 ;
    END
  END WL184
  PIN WL185
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1683.550 -1.950 1683.750 ;
        RECT -3.750 1682.950 -1.750 1683.550 ;
        RECT -3.750 1682.750 -1.950 1682.950 ;
    END
  END WL185
  PIN WL186
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1681.300 -1.950 1681.500 ;
        RECT -3.750 1680.700 -1.750 1681.300 ;
        RECT -3.750 1680.500 -1.950 1680.700 ;
    END
  END WL186
  PIN WL187
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1679.950 -1.950 1680.150 ;
        RECT -3.750 1679.350 -1.750 1679.950 ;
        RECT -3.750 1679.150 -1.950 1679.350 ;
    END
  END WL187
  PIN WL188
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1677.700 -1.950 1677.900 ;
        RECT -3.750 1677.100 -1.750 1677.700 ;
        RECT -3.750 1676.900 -1.950 1677.100 ;
    END
  END WL188
  PIN WL189
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1676.350 -1.950 1676.550 ;
        RECT -3.750 1675.750 -1.750 1676.350 ;
        RECT -3.750 1675.550 -1.950 1675.750 ;
    END
  END WL189
  PIN WL190
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1674.100 -1.950 1674.300 ;
        RECT -3.750 1673.500 -1.750 1674.100 ;
        RECT -3.750 1673.300 -1.950 1673.500 ;
    END
  END WL190
  PIN WL191
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1672.750 -1.950 1672.950 ;
        RECT -3.750 1672.150 -1.750 1672.750 ;
        RECT -3.750 1671.950 -1.950 1672.150 ;
    END
  END WL191
  PIN WL192
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1670.500 -1.950 1670.700 ;
        RECT -3.750 1669.900 -1.750 1670.500 ;
        RECT -3.750 1669.700 -1.950 1669.900 ;
    END
  END WL192
  PIN WL193
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1669.150 -1.950 1669.350 ;
        RECT -3.750 1668.550 -1.750 1669.150 ;
        RECT -3.750 1668.350 -1.950 1668.550 ;
    END
  END WL193
  PIN WL194
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1666.900 -1.950 1667.100 ;
        RECT -3.750 1666.300 -1.750 1666.900 ;
        RECT -3.750 1666.100 -1.950 1666.300 ;
    END
  END WL194
  PIN WL195
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1665.550 -1.950 1665.750 ;
        RECT -3.750 1664.950 -1.750 1665.550 ;
        RECT -3.750 1664.750 -1.950 1664.950 ;
    END
  END WL195
  PIN WL196
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1663.300 -1.950 1663.500 ;
        RECT -3.750 1662.700 -1.750 1663.300 ;
        RECT -3.750 1662.500 -1.950 1662.700 ;
    END
  END WL196
  PIN WL197
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1661.950 -1.950 1662.150 ;
        RECT -3.750 1661.350 -1.750 1661.950 ;
        RECT -3.750 1661.150 -1.950 1661.350 ;
    END
  END WL197
  PIN WL198
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1659.700 -1.950 1659.900 ;
        RECT -3.750 1659.100 -1.750 1659.700 ;
        RECT -3.750 1658.900 -1.950 1659.100 ;
    END
  END WL198
  PIN WL199
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1658.350 -1.950 1658.550 ;
        RECT -3.750 1657.750 -1.750 1658.350 ;
        RECT -3.750 1657.550 -1.950 1657.750 ;
    END
  END WL199
  PIN WL200
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1656.100 -1.950 1656.300 ;
        RECT -3.750 1655.500 -1.750 1656.100 ;
        RECT -3.750 1655.300 -1.950 1655.500 ;
    END
  END WL200
  PIN WL201
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1654.750 -1.950 1654.950 ;
        RECT -3.750 1654.150 -1.750 1654.750 ;
        RECT -3.750 1653.950 -1.950 1654.150 ;
    END
  END WL201
  PIN WL202
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1652.500 -1.950 1652.700 ;
        RECT -3.750 1651.900 -1.750 1652.500 ;
        RECT -3.750 1651.700 -1.950 1651.900 ;
    END
  END WL202
  PIN WL203
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1651.150 -1.950 1651.350 ;
        RECT -3.750 1650.550 -1.750 1651.150 ;
        RECT -3.750 1650.350 -1.950 1650.550 ;
    END
  END WL203
  PIN WL204
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1648.900 -1.950 1649.100 ;
        RECT -3.750 1648.300 -1.750 1648.900 ;
        RECT -3.750 1648.100 -1.950 1648.300 ;
    END
  END WL204
  PIN WL205
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1647.550 -1.950 1647.750 ;
        RECT -3.750 1646.950 -1.750 1647.550 ;
        RECT -3.750 1646.750 -1.950 1646.950 ;
    END
  END WL205
  PIN WL206
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1645.300 -1.950 1645.500 ;
        RECT -3.750 1644.700 -1.750 1645.300 ;
        RECT -3.750 1644.500 -1.950 1644.700 ;
    END
  END WL206
  PIN WL207
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1643.950 -1.950 1644.150 ;
        RECT -3.750 1643.350 -1.750 1643.950 ;
        RECT -3.750 1643.150 -1.950 1643.350 ;
    END
  END WL207
  PIN WL208
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1641.700 -1.950 1641.900 ;
        RECT -3.750 1641.100 -1.750 1641.700 ;
        RECT -3.750 1640.900 -1.950 1641.100 ;
    END
  END WL208
  PIN WL209
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1640.350 -1.950 1640.550 ;
        RECT -3.750 1639.750 -1.750 1640.350 ;
        RECT -3.750 1639.550 -1.950 1639.750 ;
    END
  END WL209
  PIN WL210
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1638.100 -1.950 1638.300 ;
        RECT -3.750 1637.500 -1.750 1638.100 ;
        RECT -3.750 1637.300 -1.950 1637.500 ;
    END
  END WL210
  PIN WL211
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1636.750 -1.950 1636.950 ;
        RECT -3.750 1636.150 -1.750 1636.750 ;
        RECT -3.750 1635.950 -1.950 1636.150 ;
    END
  END WL211
  PIN WL212
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1634.500 -1.950 1634.700 ;
        RECT -3.750 1633.900 -1.750 1634.500 ;
        RECT -3.750 1633.700 -1.950 1633.900 ;
    END
  END WL212
  PIN WL213
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1633.150 -1.950 1633.350 ;
        RECT -3.750 1632.550 -1.750 1633.150 ;
        RECT -3.750 1632.350 -1.950 1632.550 ;
    END
  END WL213
  PIN WL214
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1630.900 -1.950 1631.100 ;
        RECT -3.750 1630.300 -1.750 1630.900 ;
        RECT -3.750 1630.100 -1.950 1630.300 ;
    END
  END WL214
  PIN WL215
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1629.550 -1.950 1629.750 ;
        RECT -3.750 1628.950 -1.750 1629.550 ;
        RECT -3.750 1628.750 -1.950 1628.950 ;
    END
  END WL215
  PIN WL216
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1627.300 -1.950 1627.500 ;
        RECT -3.750 1626.700 -1.750 1627.300 ;
        RECT -3.750 1626.500 -1.950 1626.700 ;
    END
  END WL216
  PIN WL217
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1625.950 -1.950 1626.150 ;
        RECT -3.750 1625.350 -1.750 1625.950 ;
        RECT -3.750 1625.150 -1.950 1625.350 ;
    END
  END WL217
  PIN WL218
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1623.700 -1.950 1623.900 ;
        RECT -3.750 1623.100 -1.750 1623.700 ;
        RECT -3.750 1622.900 -1.950 1623.100 ;
    END
  END WL218
  PIN WL219
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1622.350 -1.950 1622.550 ;
        RECT -3.750 1621.750 -1.750 1622.350 ;
        RECT -3.750 1621.550 -1.950 1621.750 ;
    END
  END WL219
  PIN WL220
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1620.100 -1.950 1620.300 ;
        RECT -3.750 1619.500 -1.750 1620.100 ;
        RECT -3.750 1619.300 -1.950 1619.500 ;
    END
  END WL220
  PIN WL221
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1618.750 -1.950 1618.950 ;
        RECT -3.750 1618.150 -1.750 1618.750 ;
        RECT -3.750 1617.950 -1.950 1618.150 ;
    END
  END WL221
  PIN WL222
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1616.500 -1.950 1616.700 ;
        RECT -3.750 1615.900 -1.750 1616.500 ;
        RECT -3.750 1615.700 -1.950 1615.900 ;
    END
  END WL222
  PIN WL223
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1615.150 -1.950 1615.350 ;
        RECT -3.750 1614.550 -1.750 1615.150 ;
        RECT -3.750 1614.350 -1.950 1614.550 ;
    END
  END WL223
  PIN WL224
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1612.350 -1.950 1612.550 ;
        RECT -3.750 1611.750 -1.750 1612.350 ;
        RECT -3.750 1611.550 -1.950 1611.750 ;
    END
  END WL224
  PIN WL225
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1611.000 -1.950 1611.200 ;
        RECT -3.750 1610.400 -1.750 1611.000 ;
        RECT -3.750 1610.200 -1.950 1610.400 ;
    END
  END WL225
  PIN WL226
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1608.750 -1.950 1608.950 ;
        RECT -3.750 1608.150 -1.750 1608.750 ;
        RECT -3.750 1607.950 -1.950 1608.150 ;
    END
  END WL226
  PIN WL227
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1607.400 -1.950 1607.600 ;
        RECT -3.750 1606.800 -1.750 1607.400 ;
        RECT -3.750 1606.600 -1.950 1606.800 ;
    END
  END WL227
  PIN WL228
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1605.150 -1.950 1605.350 ;
        RECT -3.750 1604.550 -1.750 1605.150 ;
        RECT -3.750 1604.350 -1.950 1604.550 ;
    END
  END WL228
  PIN WL229
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1603.800 -1.950 1604.000 ;
        RECT -3.750 1603.200 -1.750 1603.800 ;
        RECT -3.750 1603.000 -1.950 1603.200 ;
    END
  END WL229
  PIN WL230
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1601.550 -1.950 1601.750 ;
        RECT -3.750 1600.950 -1.750 1601.550 ;
        RECT -3.750 1600.750 -1.950 1600.950 ;
    END
  END WL230
  PIN WL231
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1600.200 -1.950 1600.400 ;
        RECT -3.750 1599.600 -1.750 1600.200 ;
        RECT -3.750 1599.400 -1.950 1599.600 ;
    END
  END WL231
  PIN WL232
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1597.950 -1.950 1598.150 ;
        RECT -3.750 1597.350 -1.750 1597.950 ;
        RECT -3.750 1597.150 -1.950 1597.350 ;
    END
  END WL232
  PIN WL233
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1596.600 -1.950 1596.800 ;
        RECT -3.750 1596.000 -1.750 1596.600 ;
        RECT -3.750 1595.800 -1.950 1596.000 ;
    END
  END WL233
  PIN WL234
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1594.350 -1.950 1594.550 ;
        RECT -3.750 1593.750 -1.750 1594.350 ;
        RECT -3.750 1593.550 -1.950 1593.750 ;
    END
  END WL234
  PIN WL235
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1593.000 -1.950 1593.200 ;
        RECT -3.750 1592.400 -1.750 1593.000 ;
        RECT -3.750 1592.200 -1.950 1592.400 ;
    END
  END WL235
  PIN WL236
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1590.750 -1.950 1590.950 ;
        RECT -3.750 1590.150 -1.750 1590.750 ;
        RECT -3.750 1589.950 -1.950 1590.150 ;
    END
  END WL236
  PIN WL237
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1589.400 -1.950 1589.600 ;
        RECT -3.750 1588.800 -1.750 1589.400 ;
        RECT -3.750 1588.600 -1.950 1588.800 ;
    END
  END WL237
  PIN WL238
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1587.150 -1.950 1587.350 ;
        RECT -3.750 1586.550 -1.750 1587.150 ;
        RECT -3.750 1586.350 -1.950 1586.550 ;
    END
  END WL238
  PIN WL239
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1585.800 -1.950 1586.000 ;
        RECT -3.750 1585.200 -1.750 1585.800 ;
        RECT -3.750 1585.000 -1.950 1585.200 ;
    END
  END WL239
  PIN WL240
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1583.550 -1.950 1583.750 ;
        RECT -3.750 1582.950 -1.750 1583.550 ;
        RECT -3.750 1582.750 -1.950 1582.950 ;
    END
  END WL240
  PIN WL241
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1582.200 -1.950 1582.400 ;
        RECT -3.750 1581.600 -1.750 1582.200 ;
        RECT -3.750 1581.400 -1.950 1581.600 ;
    END
  END WL241
  PIN WL242
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1579.950 -1.950 1580.150 ;
        RECT -3.750 1579.350 -1.750 1579.950 ;
        RECT -3.750 1579.150 -1.950 1579.350 ;
    END
  END WL242
  PIN WL243
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1578.600 -1.950 1578.800 ;
        RECT -3.750 1578.000 -1.750 1578.600 ;
        RECT -3.750 1577.800 -1.950 1578.000 ;
    END
  END WL243
  PIN WL244
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1576.350 -1.950 1576.550 ;
        RECT -3.750 1575.750 -1.750 1576.350 ;
        RECT -3.750 1575.550 -1.950 1575.750 ;
    END
  END WL244
  PIN WL245
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1575.000 -1.950 1575.200 ;
        RECT -3.750 1574.400 -1.750 1575.000 ;
        RECT -3.750 1574.200 -1.950 1574.400 ;
    END
  END WL245
  PIN WL246
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1572.750 -1.950 1572.950 ;
        RECT -3.750 1572.150 -1.750 1572.750 ;
        RECT -3.750 1571.950 -1.950 1572.150 ;
    END
  END WL246
  PIN WL247
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1571.400 -1.950 1571.600 ;
        RECT -3.750 1570.800 -1.750 1571.400 ;
        RECT -3.750 1570.600 -1.950 1570.800 ;
    END
  END WL247
  PIN WL248
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1569.150 -1.950 1569.350 ;
        RECT -3.750 1568.550 -1.750 1569.150 ;
        RECT -3.750 1568.350 -1.950 1568.550 ;
    END
  END WL248
  PIN WL249
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1567.800 -1.950 1568.000 ;
        RECT -3.750 1567.200 -1.750 1567.800 ;
        RECT -3.750 1567.000 -1.950 1567.200 ;
    END
  END WL249
  PIN WL250
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1565.550 -1.950 1565.750 ;
        RECT -3.750 1564.950 -1.750 1565.550 ;
        RECT -3.750 1564.750 -1.950 1564.950 ;
    END
  END WL250
  PIN WL251
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1564.200 -1.950 1564.400 ;
        RECT -3.750 1563.600 -1.750 1564.200 ;
        RECT -3.750 1563.400 -1.950 1563.600 ;
    END
  END WL251
  PIN WL252
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1561.950 -1.950 1562.150 ;
        RECT -3.750 1561.350 -1.750 1561.950 ;
        RECT -3.750 1561.150 -1.950 1561.350 ;
    END
  END WL252
  PIN WL253
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1560.600 -1.950 1560.800 ;
        RECT -3.750 1560.000 -1.750 1560.600 ;
        RECT -3.750 1559.800 -1.950 1560.000 ;
    END
  END WL253
  PIN WL254
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1558.350 -1.950 1558.550 ;
        RECT -3.750 1557.750 -1.750 1558.350 ;
        RECT -3.750 1557.550 -1.950 1557.750 ;
    END
  END WL254
  PIN WL255
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1557.000 -1.950 1557.200 ;
        RECT -3.750 1556.400 -1.750 1557.000 ;
        RECT -3.750 1556.200 -1.950 1556.400 ;
    END
  END WL255
  PIN WL256
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1554.750 -1.950 1554.950 ;
        RECT -3.750 1554.150 -1.750 1554.750 ;
        RECT -3.750 1553.950 -1.950 1554.150 ;
    END
  END WL256
  PIN WL257
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1553.400 -1.950 1553.600 ;
        RECT -3.750 1552.800 -1.750 1553.400 ;
        RECT -3.750 1552.600 -1.950 1552.800 ;
    END
  END WL257
  PIN WL258
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1551.150 -1.950 1551.350 ;
        RECT -3.750 1550.550 -1.750 1551.150 ;
        RECT -3.750 1550.350 -1.950 1550.550 ;
    END
  END WL258
  PIN WL259
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1549.800 -1.950 1550.000 ;
        RECT -3.750 1549.200 -1.750 1549.800 ;
        RECT -3.750 1549.000 -1.950 1549.200 ;
    END
  END WL259
  PIN WL260
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1547.550 -1.950 1547.750 ;
        RECT -3.750 1546.950 -1.750 1547.550 ;
        RECT -3.750 1546.750 -1.950 1546.950 ;
    END
  END WL260
  PIN WL261
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1546.200 -1.950 1546.400 ;
        RECT -3.750 1545.600 -1.750 1546.200 ;
        RECT -3.750 1545.400 -1.950 1545.600 ;
    END
  END WL261
  PIN WL262
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1543.950 -1.950 1544.150 ;
        RECT -3.750 1543.350 -1.750 1543.950 ;
        RECT -3.750 1543.150 -1.950 1543.350 ;
    END
  END WL262
  PIN WL263
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1542.600 -1.950 1542.800 ;
        RECT -3.750 1542.000 -1.750 1542.600 ;
        RECT -3.750 1541.800 -1.950 1542.000 ;
    END
  END WL263
  PIN WL264
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1540.350 -1.950 1540.550 ;
        RECT -3.750 1539.750 -1.750 1540.350 ;
        RECT -3.750 1539.550 -1.950 1539.750 ;
    END
  END WL264
  PIN WL265
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1539.000 -1.950 1539.200 ;
        RECT -3.750 1538.400 -1.750 1539.000 ;
        RECT -3.750 1538.200 -1.950 1538.400 ;
    END
  END WL265
  PIN WL266
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1536.750 -1.950 1536.950 ;
        RECT -3.750 1536.150 -1.750 1536.750 ;
        RECT -3.750 1535.950 -1.950 1536.150 ;
    END
  END WL266
  PIN WL267
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1535.400 -1.950 1535.600 ;
        RECT -3.750 1534.800 -1.750 1535.400 ;
        RECT -3.750 1534.600 -1.950 1534.800 ;
    END
  END WL267
  PIN WL268
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1533.150 -1.950 1533.350 ;
        RECT -3.750 1532.550 -1.750 1533.150 ;
        RECT -3.750 1532.350 -1.950 1532.550 ;
    END
  END WL268
  PIN WL269
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1531.800 -1.950 1532.000 ;
        RECT -3.750 1531.200 -1.750 1531.800 ;
        RECT -3.750 1531.000 -1.950 1531.200 ;
    END
  END WL269
  PIN WL270
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1529.550 -1.950 1529.750 ;
        RECT -3.750 1528.950 -1.750 1529.550 ;
        RECT -3.750 1528.750 -1.950 1528.950 ;
    END
  END WL270
  PIN WL271
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1528.200 -1.950 1528.400 ;
        RECT -3.750 1527.600 -1.750 1528.200 ;
        RECT -3.750 1527.400 -1.950 1527.600 ;
    END
  END WL271
  PIN WL272
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1525.950 -1.950 1526.150 ;
        RECT -3.750 1525.350 -1.750 1525.950 ;
        RECT -3.750 1525.150 -1.950 1525.350 ;
    END
  END WL272
  PIN WL273
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1524.600 -1.950 1524.800 ;
        RECT -3.750 1524.000 -1.750 1524.600 ;
        RECT -3.750 1523.800 -1.950 1524.000 ;
    END
  END WL273
  PIN WL274
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1522.350 -1.950 1522.550 ;
        RECT -3.750 1521.750 -1.750 1522.350 ;
        RECT -3.750 1521.550 -1.950 1521.750 ;
    END
  END WL274
  PIN WL275
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1521.000 -1.950 1521.200 ;
        RECT -3.750 1520.400 -1.750 1521.000 ;
        RECT -3.750 1520.200 -1.950 1520.400 ;
    END
  END WL275
  PIN WL276
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1518.750 -1.950 1518.950 ;
        RECT -3.750 1518.150 -1.750 1518.750 ;
        RECT -3.750 1517.950 -1.950 1518.150 ;
    END
  END WL276
  PIN WL277
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1517.400 -1.950 1517.600 ;
        RECT -3.750 1516.800 -1.750 1517.400 ;
        RECT -3.750 1516.600 -1.950 1516.800 ;
    END
  END WL277
  PIN WL278
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1515.150 -1.950 1515.350 ;
        RECT -3.750 1514.550 -1.750 1515.150 ;
        RECT -3.750 1514.350 -1.950 1514.550 ;
    END
  END WL278
  PIN WL279
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1513.800 -1.950 1514.000 ;
        RECT -3.750 1513.200 -1.750 1513.800 ;
        RECT -3.750 1513.000 -1.950 1513.200 ;
    END
  END WL279
  PIN WL280
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1511.550 -1.950 1511.750 ;
        RECT -3.750 1510.950 -1.750 1511.550 ;
        RECT -3.750 1510.750 -1.950 1510.950 ;
    END
  END WL280
  PIN WL281
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1510.200 -1.950 1510.400 ;
        RECT -3.750 1509.600 -1.750 1510.200 ;
        RECT -3.750 1509.400 -1.950 1509.600 ;
    END
  END WL281
  PIN WL282
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1507.950 -1.950 1508.150 ;
        RECT -3.750 1507.350 -1.750 1507.950 ;
        RECT -3.750 1507.150 -1.950 1507.350 ;
    END
  END WL282
  PIN WL283
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1506.600 -1.950 1506.800 ;
        RECT -3.750 1506.000 -1.750 1506.600 ;
        RECT -3.750 1505.800 -1.950 1506.000 ;
    END
  END WL283
  PIN WL284
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1504.350 -1.950 1504.550 ;
        RECT -3.750 1503.750 -1.750 1504.350 ;
        RECT -3.750 1503.550 -1.950 1503.750 ;
    END
  END WL284
  PIN WL285
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1503.000 -1.950 1503.200 ;
        RECT -3.750 1502.400 -1.750 1503.000 ;
        RECT -3.750 1502.200 -1.950 1502.400 ;
    END
  END WL285
  PIN WL286
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1500.750 -1.950 1500.950 ;
        RECT -3.750 1500.150 -1.750 1500.750 ;
        RECT -3.750 1499.950 -1.950 1500.150 ;
    END
  END WL286
  PIN WL287
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1499.400 -1.950 1499.600 ;
        RECT -3.750 1498.800 -1.750 1499.400 ;
        RECT -3.750 1498.600 -1.950 1498.800 ;
    END
  END WL287
  PIN WL288
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1497.150 -1.950 1497.350 ;
        RECT -3.750 1496.550 -1.750 1497.150 ;
        RECT -3.750 1496.350 -1.950 1496.550 ;
    END
  END WL288
  PIN WL289
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1495.800 -1.950 1496.000 ;
        RECT -3.750 1495.200 -1.750 1495.800 ;
        RECT -3.750 1495.000 -1.950 1495.200 ;
    END
  END WL289
  PIN WL290
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1493.550 -1.950 1493.750 ;
        RECT -3.750 1492.950 -1.750 1493.550 ;
        RECT -3.750 1492.750 -1.950 1492.950 ;
    END
  END WL290
  PIN WL291
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1492.200 -1.950 1492.400 ;
        RECT -3.750 1491.600 -1.750 1492.200 ;
        RECT -3.750 1491.400 -1.950 1491.600 ;
    END
  END WL291
  PIN WL292
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1489.950 -1.950 1490.150 ;
        RECT -3.750 1489.350 -1.750 1489.950 ;
        RECT -3.750 1489.150 -1.950 1489.350 ;
    END
  END WL292
  PIN WL293
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1488.600 -1.950 1488.800 ;
        RECT -3.750 1488.000 -1.750 1488.600 ;
        RECT -3.750 1487.800 -1.950 1488.000 ;
    END
  END WL293
  PIN WL294
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1486.350 -1.950 1486.550 ;
        RECT -3.750 1485.750 -1.750 1486.350 ;
        RECT -3.750 1485.550 -1.950 1485.750 ;
    END
  END WL294
  PIN WL295
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1485.000 -1.950 1485.200 ;
        RECT -3.750 1484.400 -1.750 1485.000 ;
        RECT -3.750 1484.200 -1.950 1484.400 ;
    END
  END WL295
  PIN WL296
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1482.750 -1.950 1482.950 ;
        RECT -3.750 1482.150 -1.750 1482.750 ;
        RECT -3.750 1481.950 -1.950 1482.150 ;
    END
  END WL296
  PIN WL297
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1481.400 -1.950 1481.600 ;
        RECT -3.750 1480.800 -1.750 1481.400 ;
        RECT -3.750 1480.600 -1.950 1480.800 ;
    END
  END WL297
  PIN WL298
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1479.150 -1.950 1479.350 ;
        RECT -3.750 1478.550 -1.750 1479.150 ;
        RECT -3.750 1478.350 -1.950 1478.550 ;
    END
  END WL298
  PIN WL299
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1477.800 -1.950 1478.000 ;
        RECT -3.750 1477.200 -1.750 1477.800 ;
        RECT -3.750 1477.000 -1.950 1477.200 ;
    END
  END WL299
  PIN WL300
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1475.550 -1.950 1475.750 ;
        RECT -3.750 1474.950 -1.750 1475.550 ;
        RECT -3.750 1474.750 -1.950 1474.950 ;
    END
  END WL300
  PIN WL301
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1474.200 -1.950 1474.400 ;
        RECT -3.750 1473.600 -1.750 1474.200 ;
        RECT -3.750 1473.400 -1.950 1473.600 ;
    END
  END WL301
  PIN WL302
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1471.950 -1.950 1472.150 ;
        RECT -3.750 1471.350 -1.750 1471.950 ;
        RECT -3.750 1471.150 -1.950 1471.350 ;
    END
  END WL302
  PIN WL303
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1470.600 -1.950 1470.800 ;
        RECT -3.750 1470.000 -1.750 1470.600 ;
        RECT -3.750 1469.800 -1.950 1470.000 ;
    END
  END WL303
  PIN WL304
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1468.350 -1.950 1468.550 ;
        RECT -3.750 1467.750 -1.750 1468.350 ;
        RECT -3.750 1467.550 -1.950 1467.750 ;
    END
  END WL304
  PIN WL305
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1467.000 -1.950 1467.200 ;
        RECT -3.750 1466.400 -1.750 1467.000 ;
        RECT -3.750 1466.200 -1.950 1466.400 ;
    END
  END WL305
  PIN WL306
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1464.750 -1.950 1464.950 ;
        RECT -3.750 1464.150 -1.750 1464.750 ;
        RECT -3.750 1463.950 -1.950 1464.150 ;
    END
  END WL306
  PIN WL307
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1463.400 -1.950 1463.600 ;
        RECT -3.750 1462.800 -1.750 1463.400 ;
        RECT -3.750 1462.600 -1.950 1462.800 ;
    END
  END WL307
  PIN WL308
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1461.150 -1.950 1461.350 ;
        RECT -3.750 1460.550 -1.750 1461.150 ;
        RECT -3.750 1460.350 -1.950 1460.550 ;
    END
  END WL308
  PIN WL309
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1459.800 -1.950 1460.000 ;
        RECT -3.750 1459.200 -1.750 1459.800 ;
        RECT -3.750 1459.000 -1.950 1459.200 ;
    END
  END WL309
  PIN WL310
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1457.550 -1.950 1457.750 ;
        RECT -3.750 1456.950 -1.750 1457.550 ;
        RECT -3.750 1456.750 -1.950 1456.950 ;
    END
  END WL310
  PIN WL311
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1456.200 -1.950 1456.400 ;
        RECT -3.750 1455.600 -1.750 1456.200 ;
        RECT -3.750 1455.400 -1.950 1455.600 ;
    END
  END WL311
  PIN WL312
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1453.950 -1.950 1454.150 ;
        RECT -3.750 1453.350 -1.750 1453.950 ;
        RECT -3.750 1453.150 -1.950 1453.350 ;
    END
  END WL312
  PIN WL313
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1452.600 -1.950 1452.800 ;
        RECT -3.750 1452.000 -1.750 1452.600 ;
        RECT -3.750 1451.800 -1.950 1452.000 ;
    END
  END WL313
  PIN WL314
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1450.350 -1.950 1450.550 ;
        RECT -3.750 1449.750 -1.750 1450.350 ;
        RECT -3.750 1449.550 -1.950 1449.750 ;
    END
  END WL314
  PIN WL315
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1449.000 -1.950 1449.200 ;
        RECT -3.750 1448.400 -1.750 1449.000 ;
        RECT -3.750 1448.200 -1.950 1448.400 ;
    END
  END WL315
  PIN WL316
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1446.750 -1.950 1446.950 ;
        RECT -3.750 1446.150 -1.750 1446.750 ;
        RECT -3.750 1445.950 -1.950 1446.150 ;
    END
  END WL316
  PIN WL317
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1445.400 -1.950 1445.600 ;
        RECT -3.750 1444.800 -1.750 1445.400 ;
        RECT -3.750 1444.600 -1.950 1444.800 ;
    END
  END WL317
  PIN WL318
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1443.150 -1.950 1443.350 ;
        RECT -3.750 1442.550 -1.750 1443.150 ;
        RECT -3.750 1442.350 -1.950 1442.550 ;
    END
  END WL318
  PIN WL319
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1441.800 -1.950 1442.000 ;
        RECT -3.750 1441.200 -1.750 1441.800 ;
        RECT -3.750 1441.000 -1.950 1441.200 ;
    END
  END WL319
  PIN WL320
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1439.550 -1.950 1439.750 ;
        RECT -3.750 1438.950 -1.750 1439.550 ;
        RECT -3.750 1438.750 -1.950 1438.950 ;
    END
  END WL320
  PIN WL321
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1438.200 -1.950 1438.400 ;
        RECT -3.750 1437.600 -1.750 1438.200 ;
        RECT -3.750 1437.400 -1.950 1437.600 ;
    END
  END WL321
  PIN WL322
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1435.950 -1.950 1436.150 ;
        RECT -3.750 1435.350 -1.750 1435.950 ;
        RECT -3.750 1435.150 -1.950 1435.350 ;
    END
  END WL322
  PIN WL323
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1434.600 -1.950 1434.800 ;
        RECT -3.750 1434.000 -1.750 1434.600 ;
        RECT -3.750 1433.800 -1.950 1434.000 ;
    END
  END WL323
  PIN WL324
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1432.350 -1.950 1432.550 ;
        RECT -3.750 1431.750 -1.750 1432.350 ;
        RECT -3.750 1431.550 -1.950 1431.750 ;
    END
  END WL324
  PIN WL325
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1431.000 -1.950 1431.200 ;
        RECT -3.750 1430.400 -1.750 1431.000 ;
        RECT -3.750 1430.200 -1.950 1430.400 ;
    END
  END WL325
  PIN WL326
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1428.750 -1.950 1428.950 ;
        RECT -3.750 1428.150 -1.750 1428.750 ;
        RECT -3.750 1427.950 -1.950 1428.150 ;
    END
  END WL326
  PIN WL327
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1427.400 -1.950 1427.600 ;
        RECT -3.750 1426.800 -1.750 1427.400 ;
        RECT -3.750 1426.600 -1.950 1426.800 ;
    END
  END WL327
  PIN WL328
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1425.150 -1.950 1425.350 ;
        RECT -3.750 1424.550 -1.750 1425.150 ;
        RECT -3.750 1424.350 -1.950 1424.550 ;
    END
  END WL328
  PIN WL329
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1423.800 -1.950 1424.000 ;
        RECT -3.750 1423.200 -1.750 1423.800 ;
        RECT -3.750 1423.000 -1.950 1423.200 ;
    END
  END WL329
  PIN WL330
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1421.550 -1.950 1421.750 ;
        RECT -3.750 1420.950 -1.750 1421.550 ;
        RECT -3.750 1420.750 -1.950 1420.950 ;
    END
  END WL330
  PIN WL331
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1420.200 -1.950 1420.400 ;
        RECT -3.750 1419.600 -1.750 1420.200 ;
        RECT -3.750 1419.400 -1.950 1419.600 ;
    END
  END WL331
  PIN WL332
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1417.950 -1.950 1418.150 ;
        RECT -3.750 1417.350 -1.750 1417.950 ;
        RECT -3.750 1417.150 -1.950 1417.350 ;
    END
  END WL332
  PIN WL333
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1416.600 -1.950 1416.800 ;
        RECT -3.750 1416.000 -1.750 1416.600 ;
        RECT -3.750 1415.800 -1.950 1416.000 ;
    END
  END WL333
  PIN WL334
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1413.800 -1.950 1414.000 ;
        RECT -3.750 1413.200 -1.750 1413.800 ;
        RECT -3.750 1413.000 -1.950 1413.200 ;
    END
  END WL334
  PIN WL335
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1412.450 -1.950 1412.650 ;
        RECT -3.750 1411.850 -1.750 1412.450 ;
        RECT -3.750 1411.650 -1.950 1411.850 ;
    END
  END WL335
  PIN WL336
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1410.200 -1.950 1410.400 ;
        RECT -3.750 1409.600 -1.750 1410.200 ;
        RECT -3.750 1409.400 -1.950 1409.600 ;
    END
  END WL336
  PIN WL337
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1408.850 -1.950 1409.050 ;
        RECT -3.750 1408.250 -1.750 1408.850 ;
        RECT -3.750 1408.050 -1.950 1408.250 ;
    END
  END WL337
  PIN WL338
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1406.600 -1.950 1406.800 ;
        RECT -3.750 1406.000 -1.750 1406.600 ;
        RECT -3.750 1405.800 -1.950 1406.000 ;
    END
  END WL338
  PIN WL339
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1405.250 -1.950 1405.450 ;
        RECT -3.750 1404.650 -1.750 1405.250 ;
        RECT -3.750 1404.450 -1.950 1404.650 ;
    END
  END WL339
  PIN WL340
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1403.000 -1.950 1403.200 ;
        RECT -3.750 1402.400 -1.750 1403.000 ;
        RECT -3.750 1402.200 -1.950 1402.400 ;
    END
  END WL340
  PIN WL341
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1401.650 -1.950 1401.850 ;
        RECT -3.750 1401.050 -1.750 1401.650 ;
        RECT -3.750 1400.850 -1.950 1401.050 ;
    END
  END WL341
  PIN WL342
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1399.400 -1.950 1399.600 ;
        RECT -3.750 1398.800 -1.750 1399.400 ;
        RECT -3.750 1398.600 -1.950 1398.800 ;
    END
  END WL342
  PIN WL343
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1398.050 -1.950 1398.250 ;
        RECT -3.750 1397.450 -1.750 1398.050 ;
        RECT -3.750 1397.250 -1.950 1397.450 ;
    END
  END WL343
  PIN WL344
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1395.800 -1.950 1396.000 ;
        RECT -3.750 1395.200 -1.750 1395.800 ;
        RECT -3.750 1395.000 -1.950 1395.200 ;
    END
  END WL344
  PIN WL345
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1394.450 -1.950 1394.650 ;
        RECT -3.750 1393.850 -1.750 1394.450 ;
        RECT -3.750 1393.650 -1.950 1393.850 ;
    END
  END WL345
  PIN WL346
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1392.200 -1.950 1392.400 ;
        RECT -3.750 1391.600 -1.750 1392.200 ;
        RECT -3.750 1391.400 -1.950 1391.600 ;
    END
  END WL346
  PIN WL347
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1390.850 -1.950 1391.050 ;
        RECT -3.750 1390.250 -1.750 1390.850 ;
        RECT -3.750 1390.050 -1.950 1390.250 ;
    END
  END WL347
  PIN WL348
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1388.600 -1.950 1388.800 ;
        RECT -3.750 1388.000 -1.750 1388.600 ;
        RECT -3.750 1387.800 -1.950 1388.000 ;
    END
  END WL348
  PIN WL349
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1387.250 -1.950 1387.450 ;
        RECT -3.750 1386.650 -1.750 1387.250 ;
        RECT -3.750 1386.450 -1.950 1386.650 ;
    END
  END WL349
  PIN WL350
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1385.000 -1.950 1385.200 ;
        RECT -3.750 1384.400 -1.750 1385.000 ;
        RECT -3.750 1384.200 -1.950 1384.400 ;
    END
  END WL350
  PIN WL351
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1383.650 -1.950 1383.850 ;
        RECT -3.750 1383.050 -1.750 1383.650 ;
        RECT -3.750 1382.850 -1.950 1383.050 ;
    END
  END WL351
  PIN WL352
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1381.400 -1.950 1381.600 ;
        RECT -3.750 1380.800 -1.750 1381.400 ;
        RECT -3.750 1380.600 -1.950 1380.800 ;
    END
  END WL352
  PIN WL353
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1380.050 -1.950 1380.250 ;
        RECT -3.750 1379.450 -1.750 1380.050 ;
        RECT -3.750 1379.250 -1.950 1379.450 ;
    END
  END WL353
  PIN WL354
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1377.800 -1.950 1378.000 ;
        RECT -3.750 1377.200 -1.750 1377.800 ;
        RECT -3.750 1377.000 -1.950 1377.200 ;
    END
  END WL354
  PIN WL355
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1376.450 -1.950 1376.650 ;
        RECT -3.750 1375.850 -1.750 1376.450 ;
        RECT -3.750 1375.650 -1.950 1375.850 ;
    END
  END WL355
  PIN WL356
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1374.200 -1.950 1374.400 ;
        RECT -3.750 1373.600 -1.750 1374.200 ;
        RECT -3.750 1373.400 -1.950 1373.600 ;
    END
  END WL356
  PIN WL357
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1372.850 -1.950 1373.050 ;
        RECT -3.750 1372.250 -1.750 1372.850 ;
        RECT -3.750 1372.050 -1.950 1372.250 ;
    END
  END WL357
  PIN WL358
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1370.600 -1.950 1370.800 ;
        RECT -3.750 1370.000 -1.750 1370.600 ;
        RECT -3.750 1369.800 -1.950 1370.000 ;
    END
  END WL358
  PIN WL359
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1369.250 -1.950 1369.450 ;
        RECT -3.750 1368.650 -1.750 1369.250 ;
        RECT -3.750 1368.450 -1.950 1368.650 ;
    END
  END WL359
  PIN WL360
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1367.000 -1.950 1367.200 ;
        RECT -3.750 1366.400 -1.750 1367.000 ;
        RECT -3.750 1366.200 -1.950 1366.400 ;
    END
  END WL360
  PIN WL361
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1365.650 -1.950 1365.850 ;
        RECT -3.750 1365.050 -1.750 1365.650 ;
        RECT -3.750 1364.850 -1.950 1365.050 ;
    END
  END WL361
  PIN WL362
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1363.400 -1.950 1363.600 ;
        RECT -3.750 1362.800 -1.750 1363.400 ;
        RECT -3.750 1362.600 -1.950 1362.800 ;
    END
  END WL362
  PIN WL363
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1362.050 -1.950 1362.250 ;
        RECT -3.750 1361.450 -1.750 1362.050 ;
        RECT -3.750 1361.250 -1.950 1361.450 ;
    END
  END WL363
  PIN WL364
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1359.800 -1.950 1360.000 ;
        RECT -3.750 1359.200 -1.750 1359.800 ;
        RECT -3.750 1359.000 -1.950 1359.200 ;
    END
  END WL364
  PIN WL365
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1358.450 -1.950 1358.650 ;
        RECT -3.750 1357.850 -1.750 1358.450 ;
        RECT -3.750 1357.650 -1.950 1357.850 ;
    END
  END WL365
  PIN WL366
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1356.200 -1.950 1356.400 ;
        RECT -3.750 1355.600 -1.750 1356.200 ;
        RECT -3.750 1355.400 -1.950 1355.600 ;
    END
  END WL366
  PIN WL367
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1354.850 -1.950 1355.050 ;
        RECT -3.750 1354.250 -1.750 1354.850 ;
        RECT -3.750 1354.050 -1.950 1354.250 ;
    END
  END WL367
  PIN WL368
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1352.600 -1.950 1352.800 ;
        RECT -3.750 1352.000 -1.750 1352.600 ;
        RECT -3.750 1351.800 -1.950 1352.000 ;
    END
  END WL368
  PIN WL369
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1351.250 -1.950 1351.450 ;
        RECT -3.750 1350.650 -1.750 1351.250 ;
        RECT -3.750 1350.450 -1.950 1350.650 ;
    END
  END WL369
  PIN WL370
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1349.000 -1.950 1349.200 ;
        RECT -3.750 1348.400 -1.750 1349.000 ;
        RECT -3.750 1348.200 -1.950 1348.400 ;
    END
  END WL370
  PIN WL371
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1347.650 -1.950 1347.850 ;
        RECT -3.750 1347.050 -1.750 1347.650 ;
        RECT -3.750 1346.850 -1.950 1347.050 ;
    END
  END WL371
  PIN WL372
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1345.400 -1.950 1345.600 ;
        RECT -3.750 1344.800 -1.750 1345.400 ;
        RECT -3.750 1344.600 -1.950 1344.800 ;
    END
  END WL372
  PIN WL373
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1344.050 -1.950 1344.250 ;
        RECT -3.750 1343.450 -1.750 1344.050 ;
        RECT -3.750 1343.250 -1.950 1343.450 ;
    END
  END WL373
  PIN WL374
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1341.800 -1.950 1342.000 ;
        RECT -3.750 1341.200 -1.750 1341.800 ;
        RECT -3.750 1341.000 -1.950 1341.200 ;
    END
  END WL374
  PIN WL375
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1340.450 -1.950 1340.650 ;
        RECT -3.750 1339.850 -1.750 1340.450 ;
        RECT -3.750 1339.650 -1.950 1339.850 ;
    END
  END WL375
  PIN WL376
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1338.200 -1.950 1338.400 ;
        RECT -3.750 1337.600 -1.750 1338.200 ;
        RECT -3.750 1337.400 -1.950 1337.600 ;
    END
  END WL376
  PIN WL377
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1336.850 -1.950 1337.050 ;
        RECT -3.750 1336.250 -1.750 1336.850 ;
        RECT -3.750 1336.050 -1.950 1336.250 ;
    END
  END WL377
  PIN WL378
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1334.600 -1.950 1334.800 ;
        RECT -3.750 1334.000 -1.750 1334.600 ;
        RECT -3.750 1333.800 -1.950 1334.000 ;
    END
  END WL378
  PIN WL379
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1333.250 -1.950 1333.450 ;
        RECT -3.750 1332.650 -1.750 1333.250 ;
        RECT -3.750 1332.450 -1.950 1332.650 ;
    END
  END WL379
  PIN WL380
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1331.000 -1.950 1331.200 ;
        RECT -3.750 1330.400 -1.750 1331.000 ;
        RECT -3.750 1330.200 -1.950 1330.400 ;
    END
  END WL380
  PIN WL381
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1329.650 -1.950 1329.850 ;
        RECT -3.750 1329.050 -1.750 1329.650 ;
        RECT -3.750 1328.850 -1.950 1329.050 ;
    END
  END WL381
  PIN WL382
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1327.400 -1.950 1327.600 ;
        RECT -3.750 1326.800 -1.750 1327.400 ;
        RECT -3.750 1326.600 -1.950 1326.800 ;
    END
  END WL382
  PIN WL383
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1326.050 -1.950 1326.250 ;
        RECT -3.750 1325.450 -1.750 1326.050 ;
        RECT -3.750 1325.250 -1.950 1325.450 ;
    END
  END WL383
  PIN WL384
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1323.800 -1.950 1324.000 ;
        RECT -3.750 1323.200 -1.750 1323.800 ;
        RECT -3.750 1323.000 -1.950 1323.200 ;
    END
  END WL384
  PIN WL385
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1322.450 -1.950 1322.650 ;
        RECT -3.750 1321.850 -1.750 1322.450 ;
        RECT -3.750 1321.650 -1.950 1321.850 ;
    END
  END WL385
  PIN WL386
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1320.200 -1.950 1320.400 ;
        RECT -3.750 1319.600 -1.750 1320.200 ;
        RECT -3.750 1319.400 -1.950 1319.600 ;
    END
  END WL386
  PIN WL387
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1318.850 -1.950 1319.050 ;
        RECT -3.750 1318.250 -1.750 1318.850 ;
        RECT -3.750 1318.050 -1.950 1318.250 ;
    END
  END WL387
  PIN WL388
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1316.600 -1.950 1316.800 ;
        RECT -3.750 1316.000 -1.750 1316.600 ;
        RECT -3.750 1315.800 -1.950 1316.000 ;
    END
  END WL388
  PIN WL389
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1315.250 -1.950 1315.450 ;
        RECT -3.750 1314.650 -1.750 1315.250 ;
        RECT -3.750 1314.450 -1.950 1314.650 ;
    END
  END WL389
  PIN WL390
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1313.000 -1.950 1313.200 ;
        RECT -3.750 1312.400 -1.750 1313.000 ;
        RECT -3.750 1312.200 -1.950 1312.400 ;
    END
  END WL390
  PIN WL391
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1311.650 -1.950 1311.850 ;
        RECT -3.750 1311.050 -1.750 1311.650 ;
        RECT -3.750 1310.850 -1.950 1311.050 ;
    END
  END WL391
  PIN WL392
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1309.400 -1.950 1309.600 ;
        RECT -3.750 1308.800 -1.750 1309.400 ;
        RECT -3.750 1308.600 -1.950 1308.800 ;
    END
  END WL392
  PIN WL393
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1308.050 -1.950 1308.250 ;
        RECT -3.750 1307.450 -1.750 1308.050 ;
        RECT -3.750 1307.250 -1.950 1307.450 ;
    END
  END WL393
  PIN WL394
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1305.800 -1.950 1306.000 ;
        RECT -3.750 1305.200 -1.750 1305.800 ;
        RECT -3.750 1305.000 -1.950 1305.200 ;
    END
  END WL394
  PIN WL395
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1304.450 -1.950 1304.650 ;
        RECT -3.750 1303.850 -1.750 1304.450 ;
        RECT -3.750 1303.650 -1.950 1303.850 ;
    END
  END WL395
  PIN WL396
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1302.200 -1.950 1302.400 ;
        RECT -3.750 1301.600 -1.750 1302.200 ;
        RECT -3.750 1301.400 -1.950 1301.600 ;
    END
  END WL396
  PIN WL397
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1300.850 -1.950 1301.050 ;
        RECT -3.750 1300.250 -1.750 1300.850 ;
        RECT -3.750 1300.050 -1.950 1300.250 ;
    END
  END WL397
  PIN WL398
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1298.600 -1.950 1298.800 ;
        RECT -3.750 1298.000 -1.750 1298.600 ;
        RECT -3.750 1297.800 -1.950 1298.000 ;
    END
  END WL398
  PIN WL399
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1297.250 -1.950 1297.450 ;
        RECT -3.750 1296.650 -1.750 1297.250 ;
        RECT -3.750 1296.450 -1.950 1296.650 ;
    END
  END WL399
  PIN WL400
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1295.000 -1.950 1295.200 ;
        RECT -3.750 1294.400 -1.750 1295.000 ;
        RECT -3.750 1294.200 -1.950 1294.400 ;
    END
  END WL400
  PIN WL401
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1293.650 -1.950 1293.850 ;
        RECT -3.750 1293.050 -1.750 1293.650 ;
        RECT -3.750 1292.850 -1.950 1293.050 ;
    END
  END WL401
  PIN WL402
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1291.400 -1.950 1291.600 ;
        RECT -3.750 1290.800 -1.750 1291.400 ;
        RECT -3.750 1290.600 -1.950 1290.800 ;
    END
  END WL402
  PIN WL403
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1290.050 -1.950 1290.250 ;
        RECT -3.750 1289.450 -1.750 1290.050 ;
        RECT -3.750 1289.250 -1.950 1289.450 ;
    END
  END WL403
  PIN WL404
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1287.800 -1.950 1288.000 ;
        RECT -3.750 1287.200 -1.750 1287.800 ;
        RECT -3.750 1287.000 -1.950 1287.200 ;
    END
  END WL404
  PIN WL405
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1286.450 -1.950 1286.650 ;
        RECT -3.750 1285.850 -1.750 1286.450 ;
        RECT -3.750 1285.650 -1.950 1285.850 ;
    END
  END WL405
  PIN WL406
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1284.200 -1.950 1284.400 ;
        RECT -3.750 1283.600 -1.750 1284.200 ;
        RECT -3.750 1283.400 -1.950 1283.600 ;
    END
  END WL406
  PIN WL407
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1282.850 -1.950 1283.050 ;
        RECT -3.750 1282.250 -1.750 1282.850 ;
        RECT -3.750 1282.050 -1.950 1282.250 ;
    END
  END WL407
  PIN WL408
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1280.600 -1.950 1280.800 ;
        RECT -3.750 1280.000 -1.750 1280.600 ;
        RECT -3.750 1279.800 -1.950 1280.000 ;
    END
  END WL408
  PIN WL409
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1279.250 -1.950 1279.450 ;
        RECT -3.750 1278.650 -1.750 1279.250 ;
        RECT -3.750 1278.450 -1.950 1278.650 ;
    END
  END WL409
  PIN WL410
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1277.000 -1.950 1277.200 ;
        RECT -3.750 1276.400 -1.750 1277.000 ;
        RECT -3.750 1276.200 -1.950 1276.400 ;
    END
  END WL410
  PIN WL411
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1275.650 -1.950 1275.850 ;
        RECT -3.750 1275.050 -1.750 1275.650 ;
        RECT -3.750 1274.850 -1.950 1275.050 ;
    END
  END WL411
  PIN WL412
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1273.400 -1.950 1273.600 ;
        RECT -3.750 1272.800 -1.750 1273.400 ;
        RECT -3.750 1272.600 -1.950 1272.800 ;
    END
  END WL412
  PIN WL413
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1272.050 -1.950 1272.250 ;
        RECT -3.750 1271.450 -1.750 1272.050 ;
        RECT -3.750 1271.250 -1.950 1271.450 ;
    END
  END WL413
  PIN WL414
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1269.800 -1.950 1270.000 ;
        RECT -3.750 1269.200 -1.750 1269.800 ;
        RECT -3.750 1269.000 -1.950 1269.200 ;
    END
  END WL414
  PIN WL415
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1268.450 -1.950 1268.650 ;
        RECT -3.750 1267.850 -1.750 1268.450 ;
        RECT -3.750 1267.650 -1.950 1267.850 ;
    END
  END WL415
  PIN WL416
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1266.200 -1.950 1266.400 ;
        RECT -3.750 1265.600 -1.750 1266.200 ;
        RECT -3.750 1265.400 -1.950 1265.600 ;
    END
  END WL416
  PIN WL417
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1264.850 -1.950 1265.050 ;
        RECT -3.750 1264.250 -1.750 1264.850 ;
        RECT -3.750 1264.050 -1.950 1264.250 ;
    END
  END WL417
  PIN WL418
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1262.600 -1.950 1262.800 ;
        RECT -3.750 1262.000 -1.750 1262.600 ;
        RECT -3.750 1261.800 -1.950 1262.000 ;
    END
  END WL418
  PIN WL419
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1261.250 -1.950 1261.450 ;
        RECT -3.750 1260.650 -1.750 1261.250 ;
        RECT -3.750 1260.450 -1.950 1260.650 ;
    END
  END WL419
  PIN WL420
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1259.000 -1.950 1259.200 ;
        RECT -3.750 1258.400 -1.750 1259.000 ;
        RECT -3.750 1258.200 -1.950 1258.400 ;
    END
  END WL420
  PIN WL421
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1257.650 -1.950 1257.850 ;
        RECT -3.750 1257.050 -1.750 1257.650 ;
        RECT -3.750 1256.850 -1.950 1257.050 ;
    END
  END WL421
  PIN WL422
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1255.400 -1.950 1255.600 ;
        RECT -3.750 1254.800 -1.750 1255.400 ;
        RECT -3.750 1254.600 -1.950 1254.800 ;
    END
  END WL422
  PIN WL423
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1254.050 -1.950 1254.250 ;
        RECT -3.750 1253.450 -1.750 1254.050 ;
        RECT -3.750 1253.250 -1.950 1253.450 ;
    END
  END WL423
  PIN WL424
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1251.800 -1.950 1252.000 ;
        RECT -3.750 1251.200 -1.750 1251.800 ;
        RECT -3.750 1251.000 -1.950 1251.200 ;
    END
  END WL424
  PIN WL425
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1250.450 -1.950 1250.650 ;
        RECT -3.750 1249.850 -1.750 1250.450 ;
        RECT -3.750 1249.650 -1.950 1249.850 ;
    END
  END WL425
  PIN WL426
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1248.200 -1.950 1248.400 ;
        RECT -3.750 1247.600 -1.750 1248.200 ;
        RECT -3.750 1247.400 -1.950 1247.600 ;
    END
  END WL426
  PIN WL427
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1246.850 -1.950 1247.050 ;
        RECT -3.750 1246.250 -1.750 1246.850 ;
        RECT -3.750 1246.050 -1.950 1246.250 ;
    END
  END WL427
  PIN WL428
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1244.600 -1.950 1244.800 ;
        RECT -3.750 1244.000 -1.750 1244.600 ;
        RECT -3.750 1243.800 -1.950 1244.000 ;
    END
  END WL428
  PIN WL429
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1243.250 -1.950 1243.450 ;
        RECT -3.750 1242.650 -1.750 1243.250 ;
        RECT -3.750 1242.450 -1.950 1242.650 ;
    END
  END WL429
  PIN WL430
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1241.000 -1.950 1241.200 ;
        RECT -3.750 1240.400 -1.750 1241.000 ;
        RECT -3.750 1240.200 -1.950 1240.400 ;
    END
  END WL430
  PIN WL431
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1239.650 -1.950 1239.850 ;
        RECT -3.750 1239.050 -1.750 1239.650 ;
        RECT -3.750 1238.850 -1.950 1239.050 ;
    END
  END WL431
  PIN WL432
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1237.400 -1.950 1237.600 ;
        RECT -3.750 1236.800 -1.750 1237.400 ;
        RECT -3.750 1236.600 -1.950 1236.800 ;
    END
  END WL432
  PIN WL433
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1236.050 -1.950 1236.250 ;
        RECT -3.750 1235.450 -1.750 1236.050 ;
        RECT -3.750 1235.250 -1.950 1235.450 ;
    END
  END WL433
  PIN WL434
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1233.800 -1.950 1234.000 ;
        RECT -3.750 1233.200 -1.750 1233.800 ;
        RECT -3.750 1233.000 -1.950 1233.200 ;
    END
  END WL434
  PIN WL435
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1232.450 -1.950 1232.650 ;
        RECT -3.750 1231.850 -1.750 1232.450 ;
        RECT -3.750 1231.650 -1.950 1231.850 ;
    END
  END WL435
  PIN WL436
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1230.200 -1.950 1230.400 ;
        RECT -3.750 1229.600 -1.750 1230.200 ;
        RECT -3.750 1229.400 -1.950 1229.600 ;
    END
  END WL436
  PIN WL437
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1228.850 -1.950 1229.050 ;
        RECT -3.750 1228.250 -1.750 1228.850 ;
        RECT -3.750 1228.050 -1.950 1228.250 ;
    END
  END WL437
  PIN WL438
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1226.600 -1.950 1226.800 ;
        RECT -3.750 1226.000 -1.750 1226.600 ;
        RECT -3.750 1225.800 -1.950 1226.000 ;
    END
  END WL438
  PIN WL439
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1225.250 -1.950 1225.450 ;
        RECT -3.750 1224.650 -1.750 1225.250 ;
        RECT -3.750 1224.450 -1.950 1224.650 ;
    END
  END WL439
  PIN WL440
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1223.000 -1.950 1223.200 ;
        RECT -3.750 1222.400 -1.750 1223.000 ;
        RECT -3.750 1222.200 -1.950 1222.400 ;
    END
  END WL440
  PIN WL441
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1221.650 -1.950 1221.850 ;
        RECT -3.750 1221.050 -1.750 1221.650 ;
        RECT -3.750 1220.850 -1.950 1221.050 ;
    END
  END WL441
  PIN WL442
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1219.400 -1.950 1219.600 ;
        RECT -3.750 1218.800 -1.750 1219.400 ;
        RECT -3.750 1218.600 -1.950 1218.800 ;
    END
  END WL442
  PIN WL443
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1218.050 -1.950 1218.250 ;
        RECT -3.750 1217.450 -1.750 1218.050 ;
        RECT -3.750 1217.250 -1.950 1217.450 ;
    END
  END WL443
  PIN WL444
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1215.250 -1.950 1215.450 ;
        RECT -3.750 1214.650 -1.750 1215.250 ;
        RECT -3.750 1214.450 -1.950 1214.650 ;
    END
  END WL444
  PIN WL445
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1213.900 -1.950 1214.100 ;
        RECT -3.750 1213.300 -1.750 1213.900 ;
        RECT -3.750 1213.100 -1.950 1213.300 ;
    END
  END WL445
  PIN WL446
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1211.650 -1.950 1211.850 ;
        RECT -3.750 1211.050 -1.750 1211.650 ;
        RECT -3.750 1210.850 -1.950 1211.050 ;
    END
  END WL446
  PIN WL447
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1210.300 -1.950 1210.500 ;
        RECT -3.750 1209.700 -1.750 1210.300 ;
        RECT -3.750 1209.500 -1.950 1209.700 ;
    END
  END WL447
  PIN WL448
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1208.050 -1.950 1208.250 ;
        RECT -3.750 1207.450 -1.750 1208.050 ;
        RECT -3.750 1207.250 -1.950 1207.450 ;
    END
  END WL448
  PIN WL449
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1206.700 -1.950 1206.900 ;
        RECT -3.750 1206.100 -1.750 1206.700 ;
        RECT -3.750 1205.900 -1.950 1206.100 ;
    END
  END WL449
  PIN WL450
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1204.450 -1.950 1204.650 ;
        RECT -3.750 1203.850 -1.750 1204.450 ;
        RECT -3.750 1203.650 -1.950 1203.850 ;
    END
  END WL450
  PIN WL451
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1203.100 -1.950 1203.300 ;
        RECT -3.750 1202.500 -1.750 1203.100 ;
        RECT -3.750 1202.300 -1.950 1202.500 ;
    END
  END WL451
  PIN WL452
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1200.850 -1.950 1201.050 ;
        RECT -3.750 1200.250 -1.750 1200.850 ;
        RECT -3.750 1200.050 -1.950 1200.250 ;
    END
  END WL452
  PIN WL453
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1199.500 -1.950 1199.700 ;
        RECT -3.750 1198.900 -1.750 1199.500 ;
        RECT -3.750 1198.700 -1.950 1198.900 ;
    END
  END WL453
  PIN WL454
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1197.250 -1.950 1197.450 ;
        RECT -3.750 1196.650 -1.750 1197.250 ;
        RECT -3.750 1196.450 -1.950 1196.650 ;
    END
  END WL454
  PIN WL455
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1195.900 -1.950 1196.100 ;
        RECT -3.750 1195.300 -1.750 1195.900 ;
        RECT -3.750 1195.100 -1.950 1195.300 ;
    END
  END WL455
  PIN WL456
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1193.650 -1.950 1193.850 ;
        RECT -3.750 1193.050 -1.750 1193.650 ;
        RECT -3.750 1192.850 -1.950 1193.050 ;
    END
  END WL456
  PIN WL457
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1192.300 -1.950 1192.500 ;
        RECT -3.750 1191.700 -1.750 1192.300 ;
        RECT -3.750 1191.500 -1.950 1191.700 ;
    END
  END WL457
  PIN WL458
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1190.050 -1.950 1190.250 ;
        RECT -3.750 1189.450 -1.750 1190.050 ;
        RECT -3.750 1189.250 -1.950 1189.450 ;
    END
  END WL458
  PIN WL459
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1188.700 -1.950 1188.900 ;
        RECT -3.750 1188.100 -1.750 1188.700 ;
        RECT -3.750 1187.900 -1.950 1188.100 ;
    END
  END WL459
  PIN WL460
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1186.450 -1.950 1186.650 ;
        RECT -3.750 1185.850 -1.750 1186.450 ;
        RECT -3.750 1185.650 -1.950 1185.850 ;
    END
  END WL460
  PIN WL461
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1185.100 -1.950 1185.300 ;
        RECT -3.750 1184.500 -1.750 1185.100 ;
        RECT -3.750 1184.300 -1.950 1184.500 ;
    END
  END WL461
  PIN WL462
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1182.850 -1.950 1183.050 ;
        RECT -3.750 1182.250 -1.750 1182.850 ;
        RECT -3.750 1182.050 -1.950 1182.250 ;
    END
  END WL462
  PIN WL463
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1181.500 -1.950 1181.700 ;
        RECT -3.750 1180.900 -1.750 1181.500 ;
        RECT -3.750 1180.700 -1.950 1180.900 ;
    END
  END WL463
  PIN WL464
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1179.250 -1.950 1179.450 ;
        RECT -3.750 1178.650 -1.750 1179.250 ;
        RECT -3.750 1178.450 -1.950 1178.650 ;
    END
  END WL464
  PIN WL465
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1177.900 -1.950 1178.100 ;
        RECT -3.750 1177.300 -1.750 1177.900 ;
        RECT -3.750 1177.100 -1.950 1177.300 ;
    END
  END WL465
  PIN WL466
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1175.650 -1.950 1175.850 ;
        RECT -3.750 1175.050 -1.750 1175.650 ;
        RECT -3.750 1174.850 -1.950 1175.050 ;
    END
  END WL466
  PIN WL467
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1174.300 -1.950 1174.500 ;
        RECT -3.750 1173.700 -1.750 1174.300 ;
        RECT -3.750 1173.500 -1.950 1173.700 ;
    END
  END WL467
  PIN WL468
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1172.050 -1.950 1172.250 ;
        RECT -3.750 1171.450 -1.750 1172.050 ;
        RECT -3.750 1171.250 -1.950 1171.450 ;
    END
  END WL468
  PIN WL469
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1170.700 -1.950 1170.900 ;
        RECT -3.750 1170.100 -1.750 1170.700 ;
        RECT -3.750 1169.900 -1.950 1170.100 ;
    END
  END WL469
  PIN WL470
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1168.450 -1.950 1168.650 ;
        RECT -3.750 1167.850 -1.750 1168.450 ;
        RECT -3.750 1167.650 -1.950 1167.850 ;
    END
  END WL470
  PIN WL471
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1167.100 -1.950 1167.300 ;
        RECT -3.750 1166.500 -1.750 1167.100 ;
        RECT -3.750 1166.300 -1.950 1166.500 ;
    END
  END WL471
  PIN WL472
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1164.850 -1.950 1165.050 ;
        RECT -3.750 1164.250 -1.750 1164.850 ;
        RECT -3.750 1164.050 -1.950 1164.250 ;
    END
  END WL472
  PIN WL473
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1163.500 -1.950 1163.700 ;
        RECT -3.750 1162.900 -1.750 1163.500 ;
        RECT -3.750 1162.700 -1.950 1162.900 ;
    END
  END WL473
  PIN WL474
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1161.250 -1.950 1161.450 ;
        RECT -3.750 1160.650 -1.750 1161.250 ;
        RECT -3.750 1160.450 -1.950 1160.650 ;
    END
  END WL474
  PIN WL475
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1159.900 -1.950 1160.100 ;
        RECT -3.750 1159.300 -1.750 1159.900 ;
        RECT -3.750 1159.100 -1.950 1159.300 ;
    END
  END WL475
  PIN WL476
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1157.650 -1.950 1157.850 ;
        RECT -3.750 1157.050 -1.750 1157.650 ;
        RECT -3.750 1156.850 -1.950 1157.050 ;
    END
  END WL476
  PIN WL477
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1156.300 -1.950 1156.500 ;
        RECT -3.750 1155.700 -1.750 1156.300 ;
        RECT -3.750 1155.500 -1.950 1155.700 ;
    END
  END WL477
  PIN WL478
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1154.050 -1.950 1154.250 ;
        RECT -3.750 1153.450 -1.750 1154.050 ;
        RECT -3.750 1153.250 -1.950 1153.450 ;
    END
  END WL478
  PIN WL479
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1152.700 -1.950 1152.900 ;
        RECT -3.750 1152.100 -1.750 1152.700 ;
        RECT -3.750 1151.900 -1.950 1152.100 ;
    END
  END WL479
  PIN WL480
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1150.450 -1.950 1150.650 ;
        RECT -3.750 1149.850 -1.750 1150.450 ;
        RECT -3.750 1149.650 -1.950 1149.850 ;
    END
  END WL480
  PIN WL481
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1149.100 -1.950 1149.300 ;
        RECT -3.750 1148.500 -1.750 1149.100 ;
        RECT -3.750 1148.300 -1.950 1148.500 ;
    END
  END WL481
  PIN WL482
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1146.850 -1.950 1147.050 ;
        RECT -3.750 1146.250 -1.750 1146.850 ;
        RECT -3.750 1146.050 -1.950 1146.250 ;
    END
  END WL482
  PIN WL483
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1145.500 -1.950 1145.700 ;
        RECT -3.750 1144.900 -1.750 1145.500 ;
        RECT -3.750 1144.700 -1.950 1144.900 ;
    END
  END WL483
  PIN WL484
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1143.250 -1.950 1143.450 ;
        RECT -3.750 1142.650 -1.750 1143.250 ;
        RECT -3.750 1142.450 -1.950 1142.650 ;
    END
  END WL484
  PIN WL485
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1141.900 -1.950 1142.100 ;
        RECT -3.750 1141.300 -1.750 1141.900 ;
        RECT -3.750 1141.100 -1.950 1141.300 ;
    END
  END WL485
  PIN WL486
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1139.650 -1.950 1139.850 ;
        RECT -3.750 1139.050 -1.750 1139.650 ;
        RECT -3.750 1138.850 -1.950 1139.050 ;
    END
  END WL486
  PIN WL487
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1138.300 -1.950 1138.500 ;
        RECT -3.750 1137.700 -1.750 1138.300 ;
        RECT -3.750 1137.500 -1.950 1137.700 ;
    END
  END WL487
  PIN WL488
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1136.050 -1.950 1136.250 ;
        RECT -3.750 1135.450 -1.750 1136.050 ;
        RECT -3.750 1135.250 -1.950 1135.450 ;
    END
  END WL488
  PIN WL489
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1134.700 -1.950 1134.900 ;
        RECT -3.750 1134.100 -1.750 1134.700 ;
        RECT -3.750 1133.900 -1.950 1134.100 ;
    END
  END WL489
  PIN WL490
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1132.450 -1.950 1132.650 ;
        RECT -3.750 1131.850 -1.750 1132.450 ;
        RECT -3.750 1131.650 -1.950 1131.850 ;
    END
  END WL490
  PIN WL491
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1131.100 -1.950 1131.300 ;
        RECT -3.750 1130.500 -1.750 1131.100 ;
        RECT -3.750 1130.300 -1.950 1130.500 ;
    END
  END WL491
  PIN WL492
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1128.850 -1.950 1129.050 ;
        RECT -3.750 1128.250 -1.750 1128.850 ;
        RECT -3.750 1128.050 -1.950 1128.250 ;
    END
  END WL492
  PIN WL493
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1127.500 -1.950 1127.700 ;
        RECT -3.750 1126.900 -1.750 1127.500 ;
        RECT -3.750 1126.700 -1.950 1126.900 ;
    END
  END WL493
  PIN WL494
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1125.250 -1.950 1125.450 ;
        RECT -3.750 1124.650 -1.750 1125.250 ;
        RECT -3.750 1124.450 -1.950 1124.650 ;
    END
  END WL494
  PIN WL495
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1123.900 -1.950 1124.100 ;
        RECT -3.750 1123.300 -1.750 1123.900 ;
        RECT -3.750 1123.100 -1.950 1123.300 ;
    END
  END WL495
  PIN WL496
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1121.650 -1.950 1121.850 ;
        RECT -3.750 1121.050 -1.750 1121.650 ;
        RECT -3.750 1120.850 -1.950 1121.050 ;
    END
  END WL496
  PIN WL497
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1120.300 -1.950 1120.500 ;
        RECT -3.750 1119.700 -1.750 1120.300 ;
        RECT -3.750 1119.500 -1.950 1119.700 ;
    END
  END WL497
  PIN WL498
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1118.050 -1.950 1118.250 ;
        RECT -3.750 1117.450 -1.750 1118.050 ;
        RECT -3.750 1117.250 -1.950 1117.450 ;
    END
  END WL498
  PIN WL499
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1116.700 -1.950 1116.900 ;
        RECT -3.750 1116.100 -1.750 1116.700 ;
        RECT -3.750 1115.900 -1.950 1116.100 ;
    END
  END WL499
  PIN WL500
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1114.450 -1.950 1114.650 ;
        RECT -3.750 1113.850 -1.750 1114.450 ;
        RECT -3.750 1113.650 -1.950 1113.850 ;
    END
  END WL500
  PIN WL501
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1113.100 -1.950 1113.300 ;
        RECT -3.750 1112.500 -1.750 1113.100 ;
        RECT -3.750 1112.300 -1.950 1112.500 ;
    END
  END WL501
  PIN WL502
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1110.850 -1.950 1111.050 ;
        RECT -3.750 1110.250 -1.750 1110.850 ;
        RECT -3.750 1110.050 -1.950 1110.250 ;
    END
  END WL502
  PIN WL503
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1109.500 -1.950 1109.700 ;
        RECT -3.750 1108.900 -1.750 1109.500 ;
        RECT -3.750 1108.700 -1.950 1108.900 ;
    END
  END WL503
  PIN WL504
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1107.250 -1.950 1107.450 ;
        RECT -3.750 1106.650 -1.750 1107.250 ;
        RECT -3.750 1106.450 -1.950 1106.650 ;
    END
  END WL504
  PIN WL505
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1105.900 -1.950 1106.100 ;
        RECT -3.750 1105.300 -1.750 1105.900 ;
        RECT -3.750 1105.100 -1.950 1105.300 ;
    END
  END WL505
  PIN WL506
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1103.650 -1.950 1103.850 ;
        RECT -3.750 1103.050 -1.750 1103.650 ;
        RECT -3.750 1102.850 -1.950 1103.050 ;
    END
  END WL506
  PIN WL507
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1102.300 -1.950 1102.500 ;
        RECT -3.750 1101.700 -1.750 1102.300 ;
        RECT -3.750 1101.500 -1.950 1101.700 ;
    END
  END WL507
  PIN WL508
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1100.050 -1.950 1100.250 ;
        RECT -3.750 1099.450 -1.750 1100.050 ;
        RECT -3.750 1099.250 -1.950 1099.450 ;
    END
  END WL508
  PIN WL509
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1098.700 -1.950 1098.900 ;
        RECT -3.750 1098.100 -1.750 1098.700 ;
        RECT -3.750 1097.900 -1.950 1098.100 ;
    END
  END WL509
  PIN WL510
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1096.450 -1.950 1096.650 ;
        RECT -3.750 1095.850 -1.750 1096.450 ;
        RECT -3.750 1095.650 -1.950 1095.850 ;
    END
  END WL510
  PIN WL511
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1095.100 -1.950 1095.300 ;
        RECT -3.750 1094.500 -1.750 1095.100 ;
        RECT -3.750 1094.300 -1.950 1094.500 ;
    END
  END WL511
  PIN WL512
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1092.850 -1.950 1093.050 ;
        RECT -3.750 1092.250 -1.750 1092.850 ;
        RECT -3.750 1092.050 -1.950 1092.250 ;
    END
  END WL512
  PIN WL513
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1091.500 -1.950 1091.700 ;
        RECT -3.750 1090.900 -1.750 1091.500 ;
        RECT -3.750 1090.700 -1.950 1090.900 ;
    END
  END WL513
  PIN WL514
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1089.250 -1.950 1089.450 ;
        RECT -3.750 1088.650 -1.750 1089.250 ;
        RECT -3.750 1088.450 -1.950 1088.650 ;
    END
  END WL514
  PIN WL515
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1087.900 -1.950 1088.100 ;
        RECT -3.750 1087.300 -1.750 1087.900 ;
        RECT -3.750 1087.100 -1.950 1087.300 ;
    END
  END WL515
  PIN WL516
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1085.650 -1.950 1085.850 ;
        RECT -3.750 1085.050 -1.750 1085.650 ;
        RECT -3.750 1084.850 -1.950 1085.050 ;
    END
  END WL516
  PIN WL517
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1084.300 -1.950 1084.500 ;
        RECT -3.750 1083.700 -1.750 1084.300 ;
        RECT -3.750 1083.500 -1.950 1083.700 ;
    END
  END WL517
  PIN WL518
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1082.050 -1.950 1082.250 ;
        RECT -3.750 1081.450 -1.750 1082.050 ;
        RECT -3.750 1081.250 -1.950 1081.450 ;
    END
  END WL518
  PIN WL519
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1080.700 -1.950 1080.900 ;
        RECT -3.750 1080.100 -1.750 1080.700 ;
        RECT -3.750 1079.900 -1.950 1080.100 ;
    END
  END WL519
  PIN WL520
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1078.450 -1.950 1078.650 ;
        RECT -3.750 1077.850 -1.750 1078.450 ;
        RECT -3.750 1077.650 -1.950 1077.850 ;
    END
  END WL520
  PIN WL521
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1077.100 -1.950 1077.300 ;
        RECT -3.750 1076.500 -1.750 1077.100 ;
        RECT -3.750 1076.300 -1.950 1076.500 ;
    END
  END WL521
  PIN WL522
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1074.850 -1.950 1075.050 ;
        RECT -3.750 1074.250 -1.750 1074.850 ;
        RECT -3.750 1074.050 -1.950 1074.250 ;
    END
  END WL522
  PIN WL523
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1073.500 -1.950 1073.700 ;
        RECT -3.750 1072.900 -1.750 1073.500 ;
        RECT -3.750 1072.700 -1.950 1072.900 ;
    END
  END WL523
  PIN WL524
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1071.250 -1.950 1071.450 ;
        RECT -3.750 1070.650 -1.750 1071.250 ;
        RECT -3.750 1070.450 -1.950 1070.650 ;
    END
  END WL524
  PIN WL525
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1069.900 -1.950 1070.100 ;
        RECT -3.750 1069.300 -1.750 1069.900 ;
        RECT -3.750 1069.100 -1.950 1069.300 ;
    END
  END WL525
  PIN WL526
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1067.650 -1.950 1067.850 ;
        RECT -3.750 1067.050 -1.750 1067.650 ;
        RECT -3.750 1066.850 -1.950 1067.050 ;
    END
  END WL526
  PIN WL527
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1066.300 -1.950 1066.500 ;
        RECT -3.750 1065.700 -1.750 1066.300 ;
        RECT -3.750 1065.500 -1.950 1065.700 ;
    END
  END WL527
  PIN WL528
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1064.050 -1.950 1064.250 ;
        RECT -3.750 1063.450 -1.750 1064.050 ;
        RECT -3.750 1063.250 -1.950 1063.450 ;
    END
  END WL528
  PIN WL529
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1062.700 -1.950 1062.900 ;
        RECT -3.750 1062.100 -1.750 1062.700 ;
        RECT -3.750 1061.900 -1.950 1062.100 ;
    END
  END WL529
  PIN WL530
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1060.450 -1.950 1060.650 ;
        RECT -3.750 1059.850 -1.750 1060.450 ;
        RECT -3.750 1059.650 -1.950 1059.850 ;
    END
  END WL530
  PIN WL531
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1059.100 -1.950 1059.300 ;
        RECT -3.750 1058.500 -1.750 1059.100 ;
        RECT -3.750 1058.300 -1.950 1058.500 ;
    END
  END WL531
  PIN WL532
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1056.850 -1.950 1057.050 ;
        RECT -3.750 1056.250 -1.750 1056.850 ;
        RECT -3.750 1056.050 -1.950 1056.250 ;
    END
  END WL532
  PIN WL533
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1055.500 -1.950 1055.700 ;
        RECT -3.750 1054.900 -1.750 1055.500 ;
        RECT -3.750 1054.700 -1.950 1054.900 ;
    END
  END WL533
  PIN WL534
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1053.250 -1.950 1053.450 ;
        RECT -3.750 1052.650 -1.750 1053.250 ;
        RECT -3.750 1052.450 -1.950 1052.650 ;
    END
  END WL534
  PIN WL535
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1051.900 -1.950 1052.100 ;
        RECT -3.750 1051.300 -1.750 1051.900 ;
        RECT -3.750 1051.100 -1.950 1051.300 ;
    END
  END WL535
  PIN WL536
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1049.650 -1.950 1049.850 ;
        RECT -3.750 1049.050 -1.750 1049.650 ;
        RECT -3.750 1048.850 -1.950 1049.050 ;
    END
  END WL536
  PIN WL537
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1048.300 -1.950 1048.500 ;
        RECT -3.750 1047.700 -1.750 1048.300 ;
        RECT -3.750 1047.500 -1.950 1047.700 ;
    END
  END WL537
  PIN WL538
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1046.050 -1.950 1046.250 ;
        RECT -3.750 1045.450 -1.750 1046.050 ;
        RECT -3.750 1045.250 -1.950 1045.450 ;
    END
  END WL538
  PIN WL539
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1044.700 -1.950 1044.900 ;
        RECT -3.750 1044.100 -1.750 1044.700 ;
        RECT -3.750 1043.900 -1.950 1044.100 ;
    END
  END WL539
  PIN WL540
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1042.450 -1.950 1042.650 ;
        RECT -3.750 1041.850 -1.750 1042.450 ;
        RECT -3.750 1041.650 -1.950 1041.850 ;
    END
  END WL540
  PIN WL541
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1041.100 -1.950 1041.300 ;
        RECT -3.750 1040.500 -1.750 1041.100 ;
        RECT -3.750 1040.300 -1.950 1040.500 ;
    END
  END WL541
  PIN WL542
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1038.850 -1.950 1039.050 ;
        RECT -3.750 1038.250 -1.750 1038.850 ;
        RECT -3.750 1038.050 -1.950 1038.250 ;
    END
  END WL542
  PIN WL543
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1037.500 -1.950 1037.700 ;
        RECT -3.750 1036.900 -1.750 1037.500 ;
        RECT -3.750 1036.700 -1.950 1036.900 ;
    END
  END WL543
  PIN WL544
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1035.250 -1.950 1035.450 ;
        RECT -3.750 1034.650 -1.750 1035.250 ;
        RECT -3.750 1034.450 -1.950 1034.650 ;
    END
  END WL544
  PIN WL545
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1033.900 -1.950 1034.100 ;
        RECT -3.750 1033.300 -1.750 1033.900 ;
        RECT -3.750 1033.100 -1.950 1033.300 ;
    END
  END WL545
  PIN WL546
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1031.650 -1.950 1031.850 ;
        RECT -3.750 1031.050 -1.750 1031.650 ;
        RECT -3.750 1030.850 -1.950 1031.050 ;
    END
  END WL546
  PIN WL547
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1030.300 -1.950 1030.500 ;
        RECT -3.750 1029.700 -1.750 1030.300 ;
        RECT -3.750 1029.500 -1.950 1029.700 ;
    END
  END WL547
  PIN WL548
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1028.050 -1.950 1028.250 ;
        RECT -3.750 1027.450 -1.750 1028.050 ;
        RECT -3.750 1027.250 -1.950 1027.450 ;
    END
  END WL548
  PIN WL549
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1026.700 -1.950 1026.900 ;
        RECT -3.750 1026.100 -1.750 1026.700 ;
        RECT -3.750 1025.900 -1.950 1026.100 ;
    END
  END WL549
  PIN WL550
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1024.450 -1.950 1024.650 ;
        RECT -3.750 1023.850 -1.750 1024.450 ;
        RECT -3.750 1023.650 -1.950 1023.850 ;
    END
  END WL550
  PIN WL551
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1023.100 -1.950 1023.300 ;
        RECT -3.750 1022.500 -1.750 1023.100 ;
        RECT -3.750 1022.300 -1.950 1022.500 ;
    END
  END WL551
  PIN WL552
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1020.850 -1.950 1021.050 ;
        RECT -3.750 1020.250 -1.750 1020.850 ;
        RECT -3.750 1020.050 -1.950 1020.250 ;
    END
  END WL552
  PIN WL553
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1019.500 -1.950 1019.700 ;
        RECT -3.750 1018.900 -1.750 1019.500 ;
        RECT -3.750 1018.700 -1.950 1018.900 ;
    END
  END WL553
  PIN WL554
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1016.700 -1.950 1016.900 ;
        RECT -3.750 1016.100 -1.750 1016.700 ;
        RECT -3.750 1015.900 -1.950 1016.100 ;
    END
  END WL554
  PIN WL555
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1015.350 -1.950 1015.550 ;
        RECT -3.750 1014.750 -1.750 1015.350 ;
        RECT -3.750 1014.550 -1.950 1014.750 ;
    END
  END WL555
  PIN WL556
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1013.100 -1.950 1013.300 ;
        RECT -3.750 1012.500 -1.750 1013.100 ;
        RECT -3.750 1012.300 -1.950 1012.500 ;
    END
  END WL556
  PIN WL557
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1011.750 -1.950 1011.950 ;
        RECT -3.750 1011.150 -1.750 1011.750 ;
        RECT -3.750 1010.950 -1.950 1011.150 ;
    END
  END WL557
  PIN WL558
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1009.500 -1.950 1009.700 ;
        RECT -3.750 1008.900 -1.750 1009.500 ;
        RECT -3.750 1008.700 -1.950 1008.900 ;
    END
  END WL558
  PIN WL559
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1008.150 -1.950 1008.350 ;
        RECT -3.750 1007.550 -1.750 1008.150 ;
        RECT -3.750 1007.350 -1.950 1007.550 ;
    END
  END WL559
  PIN WL560
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1005.900 -1.950 1006.100 ;
        RECT -3.750 1005.300 -1.750 1005.900 ;
        RECT -3.750 1005.100 -1.950 1005.300 ;
    END
  END WL560
  PIN WL561
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1004.550 -1.950 1004.750 ;
        RECT -3.750 1003.950 -1.750 1004.550 ;
        RECT -3.750 1003.750 -1.950 1003.950 ;
    END
  END WL561
  PIN WL562
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1002.300 -1.950 1002.500 ;
        RECT -3.750 1001.700 -1.750 1002.300 ;
        RECT -3.750 1001.500 -1.950 1001.700 ;
    END
  END WL562
  PIN WL563
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 1000.950 -1.950 1001.150 ;
        RECT -3.750 1000.350 -1.750 1000.950 ;
        RECT -3.750 1000.150 -1.950 1000.350 ;
    END
  END WL563
  PIN WL564
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 998.700 -1.950 998.900 ;
        RECT -3.750 998.100 -1.750 998.700 ;
        RECT -3.750 997.900 -1.950 998.100 ;
    END
  END WL564
  PIN WL565
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 997.350 -1.950 997.550 ;
        RECT -3.750 996.750 -1.750 997.350 ;
        RECT -3.750 996.550 -1.950 996.750 ;
    END
  END WL565
  PIN WL566
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 995.100 -1.950 995.300 ;
        RECT -3.750 994.500 -1.750 995.100 ;
        RECT -3.750 994.300 -1.950 994.500 ;
    END
  END WL566
  PIN WL567
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 993.750 -1.950 993.950 ;
        RECT -3.750 993.150 -1.750 993.750 ;
        RECT -3.750 992.950 -1.950 993.150 ;
    END
  END WL567
  PIN WL568
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 991.500 -1.950 991.700 ;
        RECT -3.750 990.900 -1.750 991.500 ;
        RECT -3.750 990.700 -1.950 990.900 ;
    END
  END WL568
  PIN WL569
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 990.150 -1.950 990.350 ;
        RECT -3.750 989.550 -1.750 990.150 ;
        RECT -3.750 989.350 -1.950 989.550 ;
    END
  END WL569
  PIN WL570
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 987.900 -1.950 988.100 ;
        RECT -3.750 987.300 -1.750 987.900 ;
        RECT -3.750 987.100 -1.950 987.300 ;
    END
  END WL570
  PIN WL571
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 986.550 -1.950 986.750 ;
        RECT -3.750 985.950 -1.750 986.550 ;
        RECT -3.750 985.750 -1.950 985.950 ;
    END
  END WL571
  PIN WL572
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 984.300 -1.950 984.500 ;
        RECT -3.750 983.700 -1.750 984.300 ;
        RECT -3.750 983.500 -1.950 983.700 ;
    END
  END WL572
  PIN WL573
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 982.950 -1.950 983.150 ;
        RECT -3.750 982.350 -1.750 982.950 ;
        RECT -3.750 982.150 -1.950 982.350 ;
    END
  END WL573
  PIN WL574
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 980.700 -1.950 980.900 ;
        RECT -3.750 980.100 -1.750 980.700 ;
        RECT -3.750 979.900 -1.950 980.100 ;
    END
  END WL574
  PIN WL575
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 979.350 -1.950 979.550 ;
        RECT -3.750 978.750 -1.750 979.350 ;
        RECT -3.750 978.550 -1.950 978.750 ;
    END
  END WL575
  PIN WL576
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 977.100 -1.950 977.300 ;
        RECT -3.750 976.500 -1.750 977.100 ;
        RECT -3.750 976.300 -1.950 976.500 ;
    END
  END WL576
  PIN WL577
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 975.750 -1.950 975.950 ;
        RECT -3.750 975.150 -1.750 975.750 ;
        RECT -3.750 974.950 -1.950 975.150 ;
    END
  END WL577
  PIN WL578
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 973.500 -1.950 973.700 ;
        RECT -3.750 972.900 -1.750 973.500 ;
        RECT -3.750 972.700 -1.950 972.900 ;
    END
  END WL578
  PIN WL579
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 972.150 -1.950 972.350 ;
        RECT -3.750 971.550 -1.750 972.150 ;
        RECT -3.750 971.350 -1.950 971.550 ;
    END
  END WL579
  PIN WL580
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 969.900 -1.950 970.100 ;
        RECT -3.750 969.300 -1.750 969.900 ;
        RECT -3.750 969.100 -1.950 969.300 ;
    END
  END WL580
  PIN WL581
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 968.550 -1.950 968.750 ;
        RECT -3.750 967.950 -1.750 968.550 ;
        RECT -3.750 967.750 -1.950 967.950 ;
    END
  END WL581
  PIN WL582
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 966.300 -1.950 966.500 ;
        RECT -3.750 965.700 -1.750 966.300 ;
        RECT -3.750 965.500 -1.950 965.700 ;
    END
  END WL582
  PIN WL583
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 964.950 -1.950 965.150 ;
        RECT -3.750 964.350 -1.750 964.950 ;
        RECT -3.750 964.150 -1.950 964.350 ;
    END
  END WL583
  PIN WL584
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 962.700 -1.950 962.900 ;
        RECT -3.750 962.100 -1.750 962.700 ;
        RECT -3.750 961.900 -1.950 962.100 ;
    END
  END WL584
  PIN WL585
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 961.350 -1.950 961.550 ;
        RECT -3.750 960.750 -1.750 961.350 ;
        RECT -3.750 960.550 -1.950 960.750 ;
    END
  END WL585
  PIN WL586
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 959.100 -1.950 959.300 ;
        RECT -3.750 958.500 -1.750 959.100 ;
        RECT -3.750 958.300 -1.950 958.500 ;
    END
  END WL586
  PIN WL587
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 957.750 -1.950 957.950 ;
        RECT -3.750 957.150 -1.750 957.750 ;
        RECT -3.750 956.950 -1.950 957.150 ;
    END
  END WL587
  PIN WL588
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 955.500 -1.950 955.700 ;
        RECT -3.750 954.900 -1.750 955.500 ;
        RECT -3.750 954.700 -1.950 954.900 ;
    END
  END WL588
  PIN WL589
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 954.150 -1.950 954.350 ;
        RECT -3.750 953.550 -1.750 954.150 ;
        RECT -3.750 953.350 -1.950 953.550 ;
    END
  END WL589
  PIN WL590
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 951.900 -1.950 952.100 ;
        RECT -3.750 951.300 -1.750 951.900 ;
        RECT -3.750 951.100 -1.950 951.300 ;
    END
  END WL590
  PIN WL591
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 950.550 -1.950 950.750 ;
        RECT -3.750 949.950 -1.750 950.550 ;
        RECT -3.750 949.750 -1.950 949.950 ;
    END
  END WL591
  PIN WL592
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 948.300 -1.950 948.500 ;
        RECT -3.750 947.700 -1.750 948.300 ;
        RECT -3.750 947.500 -1.950 947.700 ;
    END
  END WL592
  PIN WL593
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 946.950 -1.950 947.150 ;
        RECT -3.750 946.350 -1.750 946.950 ;
        RECT -3.750 946.150 -1.950 946.350 ;
    END
  END WL593
  PIN WL594
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 944.700 -1.950 944.900 ;
        RECT -3.750 944.100 -1.750 944.700 ;
        RECT -3.750 943.900 -1.950 944.100 ;
    END
  END WL594
  PIN WL595
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 943.350 -1.950 943.550 ;
        RECT -3.750 942.750 -1.750 943.350 ;
        RECT -3.750 942.550 -1.950 942.750 ;
    END
  END WL595
  PIN WL596
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 941.100 -1.950 941.300 ;
        RECT -3.750 940.500 -1.750 941.100 ;
        RECT -3.750 940.300 -1.950 940.500 ;
    END
  END WL596
  PIN WL597
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 939.750 -1.950 939.950 ;
        RECT -3.750 939.150 -1.750 939.750 ;
        RECT -3.750 938.950 -1.950 939.150 ;
    END
  END WL597
  PIN WL598
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 937.500 -1.950 937.700 ;
        RECT -3.750 936.900 -1.750 937.500 ;
        RECT -3.750 936.700 -1.950 936.900 ;
    END
  END WL598
  PIN WL599
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 936.150 -1.950 936.350 ;
        RECT -3.750 935.550 -1.750 936.150 ;
        RECT -3.750 935.350 -1.950 935.550 ;
    END
  END WL599
  PIN WL600
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 933.900 -1.950 934.100 ;
        RECT -3.750 933.300 -1.750 933.900 ;
        RECT -3.750 933.100 -1.950 933.300 ;
    END
  END WL600
  PIN WL601
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 932.550 -1.950 932.750 ;
        RECT -3.750 931.950 -1.750 932.550 ;
        RECT -3.750 931.750 -1.950 931.950 ;
    END
  END WL601
  PIN WL602
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 930.300 -1.950 930.500 ;
        RECT -3.750 929.700 -1.750 930.300 ;
        RECT -3.750 929.500 -1.950 929.700 ;
    END
  END WL602
  PIN WL603
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 928.950 -1.950 929.150 ;
        RECT -3.750 928.350 -1.750 928.950 ;
        RECT -3.750 928.150 -1.950 928.350 ;
    END
  END WL603
  PIN WL604
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 926.700 -1.950 926.900 ;
        RECT -3.750 926.100 -1.750 926.700 ;
        RECT -3.750 925.900 -1.950 926.100 ;
    END
  END WL604
  PIN WL605
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 925.350 -1.950 925.550 ;
        RECT -3.750 924.750 -1.750 925.350 ;
        RECT -3.750 924.550 -1.950 924.750 ;
    END
  END WL605
  PIN WL606
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 923.100 -1.950 923.300 ;
        RECT -3.750 922.500 -1.750 923.100 ;
        RECT -3.750 922.300 -1.950 922.500 ;
    END
  END WL606
  PIN WL607
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 921.750 -1.950 921.950 ;
        RECT -3.750 921.150 -1.750 921.750 ;
        RECT -3.750 920.950 -1.950 921.150 ;
    END
  END WL607
  PIN WL608
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 919.500 -1.950 919.700 ;
        RECT -3.750 918.900 -1.750 919.500 ;
        RECT -3.750 918.700 -1.950 918.900 ;
    END
  END WL608
  PIN WL609
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 918.150 -1.950 918.350 ;
        RECT -3.750 917.550 -1.750 918.150 ;
        RECT -3.750 917.350 -1.950 917.550 ;
    END
  END WL609
  PIN WL610
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 915.900 -1.950 916.100 ;
        RECT -3.750 915.300 -1.750 915.900 ;
        RECT -3.750 915.100 -1.950 915.300 ;
    END
  END WL610
  PIN WL611
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 914.550 -1.950 914.750 ;
        RECT -3.750 913.950 -1.750 914.550 ;
        RECT -3.750 913.750 -1.950 913.950 ;
    END
  END WL611
  PIN WL612
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 912.300 -1.950 912.500 ;
        RECT -3.750 911.700 -1.750 912.300 ;
        RECT -3.750 911.500 -1.950 911.700 ;
    END
  END WL612
  PIN WL613
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 910.950 -1.950 911.150 ;
        RECT -3.750 910.350 -1.750 910.950 ;
        RECT -3.750 910.150 -1.950 910.350 ;
    END
  END WL613
  PIN WL614
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 908.700 -1.950 908.900 ;
        RECT -3.750 908.100 -1.750 908.700 ;
        RECT -3.750 907.900 -1.950 908.100 ;
    END
  END WL614
  PIN WL615
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 907.350 -1.950 907.550 ;
        RECT -3.750 906.750 -1.750 907.350 ;
        RECT -3.750 906.550 -1.950 906.750 ;
    END
  END WL615
  PIN WL616
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 905.100 -1.950 905.300 ;
        RECT -3.750 904.500 -1.750 905.100 ;
        RECT -3.750 904.300 -1.950 904.500 ;
    END
  END WL616
  PIN WL617
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 903.750 -1.950 903.950 ;
        RECT -3.750 903.150 -1.750 903.750 ;
        RECT -3.750 902.950 -1.950 903.150 ;
    END
  END WL617
  PIN WL618
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 901.500 -1.950 901.700 ;
        RECT -3.750 900.900 -1.750 901.500 ;
        RECT -3.750 900.700 -1.950 900.900 ;
    END
  END WL618
  PIN WL619
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 900.150 -1.950 900.350 ;
        RECT -3.750 899.550 -1.750 900.150 ;
        RECT -3.750 899.350 -1.950 899.550 ;
    END
  END WL619
  PIN WL620
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 897.900 -1.950 898.100 ;
        RECT -3.750 897.300 -1.750 897.900 ;
        RECT -3.750 897.100 -1.950 897.300 ;
    END
  END WL620
  PIN WL621
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 896.550 -1.950 896.750 ;
        RECT -3.750 895.950 -1.750 896.550 ;
        RECT -3.750 895.750 -1.950 895.950 ;
    END
  END WL621
  PIN WL622
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 894.300 -1.950 894.500 ;
        RECT -3.750 893.700 -1.750 894.300 ;
        RECT -3.750 893.500 -1.950 893.700 ;
    END
  END WL622
  PIN WL623
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 892.950 -1.950 893.150 ;
        RECT -3.750 892.350 -1.750 892.950 ;
        RECT -3.750 892.150 -1.950 892.350 ;
    END
  END WL623
  PIN WL624
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 890.700 -1.950 890.900 ;
        RECT -3.750 890.100 -1.750 890.700 ;
        RECT -3.750 889.900 -1.950 890.100 ;
    END
  END WL624
  PIN WL625
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 889.350 -1.950 889.550 ;
        RECT -3.750 888.750 -1.750 889.350 ;
        RECT -3.750 888.550 -1.950 888.750 ;
    END
  END WL625
  PIN WL626
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 887.100 -1.950 887.300 ;
        RECT -3.750 886.500 -1.750 887.100 ;
        RECT -3.750 886.300 -1.950 886.500 ;
    END
  END WL626
  PIN WL627
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 885.750 -1.950 885.950 ;
        RECT -3.750 885.150 -1.750 885.750 ;
        RECT -3.750 884.950 -1.950 885.150 ;
    END
  END WL627
  PIN WL628
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 883.500 -1.950 883.700 ;
        RECT -3.750 882.900 -1.750 883.500 ;
        RECT -3.750 882.700 -1.950 882.900 ;
    END
  END WL628
  PIN WL629
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 882.150 -1.950 882.350 ;
        RECT -3.750 881.550 -1.750 882.150 ;
        RECT -3.750 881.350 -1.950 881.550 ;
    END
  END WL629
  PIN WL630
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 879.900 -1.950 880.100 ;
        RECT -3.750 879.300 -1.750 879.900 ;
        RECT -3.750 879.100 -1.950 879.300 ;
    END
  END WL630
  PIN WL631
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 878.550 -1.950 878.750 ;
        RECT -3.750 877.950 -1.750 878.550 ;
        RECT -3.750 877.750 -1.950 877.950 ;
    END
  END WL631
  PIN WL632
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 876.300 -1.950 876.500 ;
        RECT -3.750 875.700 -1.750 876.300 ;
        RECT -3.750 875.500 -1.950 875.700 ;
    END
  END WL632
  PIN WL633
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 874.950 -1.950 875.150 ;
        RECT -3.750 874.350 -1.750 874.950 ;
        RECT -3.750 874.150 -1.950 874.350 ;
    END
  END WL633
  PIN WL634
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 872.700 -1.950 872.900 ;
        RECT -3.750 872.100 -1.750 872.700 ;
        RECT -3.750 871.900 -1.950 872.100 ;
    END
  END WL634
  PIN WL635
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 871.350 -1.950 871.550 ;
        RECT -3.750 870.750 -1.750 871.350 ;
        RECT -3.750 870.550 -1.950 870.750 ;
    END
  END WL635
  PIN WL636
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 869.100 -1.950 869.300 ;
        RECT -3.750 868.500 -1.750 869.100 ;
        RECT -3.750 868.300 -1.950 868.500 ;
    END
  END WL636
  PIN WL637
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 867.750 -1.950 867.950 ;
        RECT -3.750 867.150 -1.750 867.750 ;
        RECT -3.750 866.950 -1.950 867.150 ;
    END
  END WL637
  PIN WL638
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 865.500 -1.950 865.700 ;
        RECT -3.750 864.900 -1.750 865.500 ;
        RECT -3.750 864.700 -1.950 864.900 ;
    END
  END WL638
  PIN WL639
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 864.150 -1.950 864.350 ;
        RECT -3.750 863.550 -1.750 864.150 ;
        RECT -3.750 863.350 -1.950 863.550 ;
    END
  END WL639
  PIN WL640
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 861.900 -1.950 862.100 ;
        RECT -3.750 861.300 -1.750 861.900 ;
        RECT -3.750 861.100 -1.950 861.300 ;
    END
  END WL640
  PIN WL641
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 860.550 -1.950 860.750 ;
        RECT -3.750 859.950 -1.750 860.550 ;
        RECT -3.750 859.750 -1.950 859.950 ;
    END
  END WL641
  PIN WL642
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 858.300 -1.950 858.500 ;
        RECT -3.750 857.700 -1.750 858.300 ;
        RECT -3.750 857.500 -1.950 857.700 ;
    END
  END WL642
  PIN WL643
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 856.950 -1.950 857.150 ;
        RECT -3.750 856.350 -1.750 856.950 ;
        RECT -3.750 856.150 -1.950 856.350 ;
    END
  END WL643
  PIN WL644
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 854.700 -1.950 854.900 ;
        RECT -3.750 854.100 -1.750 854.700 ;
        RECT -3.750 853.900 -1.950 854.100 ;
    END
  END WL644
  PIN WL645
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 853.350 -1.950 853.550 ;
        RECT -3.750 852.750 -1.750 853.350 ;
        RECT -3.750 852.550 -1.950 852.750 ;
    END
  END WL645
  PIN WL646
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 851.100 -1.950 851.300 ;
        RECT -3.750 850.500 -1.750 851.100 ;
        RECT -3.750 850.300 -1.950 850.500 ;
    END
  END WL646
  PIN WL647
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 849.750 -1.950 849.950 ;
        RECT -3.750 849.150 -1.750 849.750 ;
        RECT -3.750 848.950 -1.950 849.150 ;
    END
  END WL647
  PIN WL648
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 847.500 -1.950 847.700 ;
        RECT -3.750 846.900 -1.750 847.500 ;
        RECT -3.750 846.700 -1.950 846.900 ;
    END
  END WL648
  PIN WL649
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 846.150 -1.950 846.350 ;
        RECT -3.750 845.550 -1.750 846.150 ;
        RECT -3.750 845.350 -1.950 845.550 ;
    END
  END WL649
  PIN WL650
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 843.900 -1.950 844.100 ;
        RECT -3.750 843.300 -1.750 843.900 ;
        RECT -3.750 843.100 -1.950 843.300 ;
    END
  END WL650
  PIN WL651
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 842.550 -1.950 842.750 ;
        RECT -3.750 841.950 -1.750 842.550 ;
        RECT -3.750 841.750 -1.950 841.950 ;
    END
  END WL651
  PIN WL652
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 840.300 -1.950 840.500 ;
        RECT -3.750 839.700 -1.750 840.300 ;
        RECT -3.750 839.500 -1.950 839.700 ;
    END
  END WL652
  PIN WL653
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 838.950 -1.950 839.150 ;
        RECT -3.750 838.350 -1.750 838.950 ;
        RECT -3.750 838.150 -1.950 838.350 ;
    END
  END WL653
  PIN WL654
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 836.700 -1.950 836.900 ;
        RECT -3.750 836.100 -1.750 836.700 ;
        RECT -3.750 835.900 -1.950 836.100 ;
    END
  END WL654
  PIN WL655
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 835.350 -1.950 835.550 ;
        RECT -3.750 834.750 -1.750 835.350 ;
        RECT -3.750 834.550 -1.950 834.750 ;
    END
  END WL655
  PIN WL656
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 833.100 -1.950 833.300 ;
        RECT -3.750 832.500 -1.750 833.100 ;
        RECT -3.750 832.300 -1.950 832.500 ;
    END
  END WL656
  PIN WL657
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 831.750 -1.950 831.950 ;
        RECT -3.750 831.150 -1.750 831.750 ;
        RECT -3.750 830.950 -1.950 831.150 ;
    END
  END WL657
  PIN WL658
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 829.500 -1.950 829.700 ;
        RECT -3.750 828.900 -1.750 829.500 ;
        RECT -3.750 828.700 -1.950 828.900 ;
    END
  END WL658
  PIN WL659
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 828.150 -1.950 828.350 ;
        RECT -3.750 827.550 -1.750 828.150 ;
        RECT -3.750 827.350 -1.950 827.550 ;
    END
  END WL659
  PIN WL660
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 825.900 -1.950 826.100 ;
        RECT -3.750 825.300 -1.750 825.900 ;
        RECT -3.750 825.100 -1.950 825.300 ;
    END
  END WL660
  PIN WL661
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 824.550 -1.950 824.750 ;
        RECT -3.750 823.950 -1.750 824.550 ;
        RECT -3.750 823.750 -1.950 823.950 ;
    END
  END WL661
  PIN WL662
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 822.300 -1.950 822.500 ;
        RECT -3.750 821.700 -1.750 822.300 ;
        RECT -3.750 821.500 -1.950 821.700 ;
    END
  END WL662
  PIN WL663
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 820.950 -1.950 821.150 ;
        RECT -3.750 820.350 -1.750 820.950 ;
        RECT -3.750 820.150 -1.950 820.350 ;
    END
  END WL663
  PIN WL664
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 818.150 -1.950 818.350 ;
        RECT -3.750 817.550 -1.750 818.150 ;
        RECT -3.750 817.350 -1.950 817.550 ;
    END
  END WL664
  PIN WL665
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 816.800 -1.950 817.000 ;
        RECT -3.750 816.200 -1.750 816.800 ;
        RECT -3.750 816.000 -1.950 816.200 ;
    END
  END WL665
  PIN WL666
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 814.550 -1.950 814.750 ;
        RECT -3.750 813.950 -1.750 814.550 ;
        RECT -3.750 813.750 -1.950 813.950 ;
    END
  END WL666
  PIN WL667
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 813.200 -1.950 813.400 ;
        RECT -3.750 812.600 -1.750 813.200 ;
        RECT -3.750 812.400 -1.950 812.600 ;
    END
  END WL667
  PIN WL668
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 810.950 -1.950 811.150 ;
        RECT -3.750 810.350 -1.750 810.950 ;
        RECT -3.750 810.150 -1.950 810.350 ;
    END
  END WL668
  PIN WL669
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 809.600 -1.950 809.800 ;
        RECT -3.750 809.000 -1.750 809.600 ;
        RECT -3.750 808.800 -1.950 809.000 ;
    END
  END WL669
  PIN WL670
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 807.350 -1.950 807.550 ;
        RECT -3.750 806.750 -1.750 807.350 ;
        RECT -3.750 806.550 -1.950 806.750 ;
    END
  END WL670
  PIN WL671
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 806.000 -1.950 806.200 ;
        RECT -3.750 805.400 -1.750 806.000 ;
        RECT -3.750 805.200 -1.950 805.400 ;
    END
  END WL671
  PIN WL672
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 803.750 -1.950 803.950 ;
        RECT -3.750 803.150 -1.750 803.750 ;
        RECT -3.750 802.950 -1.950 803.150 ;
    END
  END WL672
  PIN WL673
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 802.400 -1.950 802.600 ;
        RECT -3.750 801.800 -1.750 802.400 ;
        RECT -3.750 801.600 -1.950 801.800 ;
    END
  END WL673
  PIN WL674
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 800.150 -1.950 800.350 ;
        RECT -3.750 799.550 -1.750 800.150 ;
        RECT -3.750 799.350 -1.950 799.550 ;
    END
  END WL674
  PIN WL675
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 798.800 -1.950 799.000 ;
        RECT -3.750 798.200 -1.750 798.800 ;
        RECT -3.750 798.000 -1.950 798.200 ;
    END
  END WL675
  PIN WL676
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 796.550 -1.950 796.750 ;
        RECT -3.750 795.950 -1.750 796.550 ;
        RECT -3.750 795.750 -1.950 795.950 ;
    END
  END WL676
  PIN WL677
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 795.200 -1.950 795.400 ;
        RECT -3.750 794.600 -1.750 795.200 ;
        RECT -3.750 794.400 -1.950 794.600 ;
    END
  END WL677
  PIN WL678
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 792.950 -1.950 793.150 ;
        RECT -3.750 792.350 -1.750 792.950 ;
        RECT -3.750 792.150 -1.950 792.350 ;
    END
  END WL678
  PIN WL679
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 791.600 -1.950 791.800 ;
        RECT -3.750 791.000 -1.750 791.600 ;
        RECT -3.750 790.800 -1.950 791.000 ;
    END
  END WL679
  PIN WL680
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 789.350 -1.950 789.550 ;
        RECT -3.750 788.750 -1.750 789.350 ;
        RECT -3.750 788.550 -1.950 788.750 ;
    END
  END WL680
  PIN WL681
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 788.000 -1.950 788.200 ;
        RECT -3.750 787.400 -1.750 788.000 ;
        RECT -3.750 787.200 -1.950 787.400 ;
    END
  END WL681
  PIN WL682
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 785.750 -1.950 785.950 ;
        RECT -3.750 785.150 -1.750 785.750 ;
        RECT -3.750 784.950 -1.950 785.150 ;
    END
  END WL682
  PIN WL683
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 784.400 -1.950 784.600 ;
        RECT -3.750 783.800 -1.750 784.400 ;
        RECT -3.750 783.600 -1.950 783.800 ;
    END
  END WL683
  PIN WL684
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 782.150 -1.950 782.350 ;
        RECT -3.750 781.550 -1.750 782.150 ;
        RECT -3.750 781.350 -1.950 781.550 ;
    END
  END WL684
  PIN WL685
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 780.800 -1.950 781.000 ;
        RECT -3.750 780.200 -1.750 780.800 ;
        RECT -3.750 780.000 -1.950 780.200 ;
    END
  END WL685
  PIN WL686
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 778.550 -1.950 778.750 ;
        RECT -3.750 777.950 -1.750 778.550 ;
        RECT -3.750 777.750 -1.950 777.950 ;
    END
  END WL686
  PIN WL687
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 777.200 -1.950 777.400 ;
        RECT -3.750 776.600 -1.750 777.200 ;
        RECT -3.750 776.400 -1.950 776.600 ;
    END
  END WL687
  PIN WL688
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 774.950 -1.950 775.150 ;
        RECT -3.750 774.350 -1.750 774.950 ;
        RECT -3.750 774.150 -1.950 774.350 ;
    END
  END WL688
  PIN WL689
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 773.600 -1.950 773.800 ;
        RECT -3.750 773.000 -1.750 773.600 ;
        RECT -3.750 772.800 -1.950 773.000 ;
    END
  END WL689
  PIN WL690
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 771.350 -1.950 771.550 ;
        RECT -3.750 770.750 -1.750 771.350 ;
        RECT -3.750 770.550 -1.950 770.750 ;
    END
  END WL690
  PIN WL691
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 770.000 -1.950 770.200 ;
        RECT -3.750 769.400 -1.750 770.000 ;
        RECT -3.750 769.200 -1.950 769.400 ;
    END
  END WL691
  PIN WL692
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 767.750 -1.950 767.950 ;
        RECT -3.750 767.150 -1.750 767.750 ;
        RECT -3.750 766.950 -1.950 767.150 ;
    END
  END WL692
  PIN WL693
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 766.400 -1.950 766.600 ;
        RECT -3.750 765.800 -1.750 766.400 ;
        RECT -3.750 765.600 -1.950 765.800 ;
    END
  END WL693
  PIN WL694
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 764.150 -1.950 764.350 ;
        RECT -3.750 763.550 -1.750 764.150 ;
        RECT -3.750 763.350 -1.950 763.550 ;
    END
  END WL694
  PIN WL695
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 762.800 -1.950 763.000 ;
        RECT -3.750 762.200 -1.750 762.800 ;
        RECT -3.750 762.000 -1.950 762.200 ;
    END
  END WL695
  PIN WL696
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 760.550 -1.950 760.750 ;
        RECT -3.750 759.950 -1.750 760.550 ;
        RECT -3.750 759.750 -1.950 759.950 ;
    END
  END WL696
  PIN WL697
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 759.200 -1.950 759.400 ;
        RECT -3.750 758.600 -1.750 759.200 ;
        RECT -3.750 758.400 -1.950 758.600 ;
    END
  END WL697
  PIN WL698
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 756.950 -1.950 757.150 ;
        RECT -3.750 756.350 -1.750 756.950 ;
        RECT -3.750 756.150 -1.950 756.350 ;
    END
  END WL698
  PIN WL699
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 755.600 -1.950 755.800 ;
        RECT -3.750 755.000 -1.750 755.600 ;
        RECT -3.750 754.800 -1.950 755.000 ;
    END
  END WL699
  PIN WL700
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 753.350 -1.950 753.550 ;
        RECT -3.750 752.750 -1.750 753.350 ;
        RECT -3.750 752.550 -1.950 752.750 ;
    END
  END WL700
  PIN WL701
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 752.000 -1.950 752.200 ;
        RECT -3.750 751.400 -1.750 752.000 ;
        RECT -3.750 751.200 -1.950 751.400 ;
    END
  END WL701
  PIN WL702
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 749.750 -1.950 749.950 ;
        RECT -3.750 749.150 -1.750 749.750 ;
        RECT -3.750 748.950 -1.950 749.150 ;
    END
  END WL702
  PIN WL703
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 748.400 -1.950 748.600 ;
        RECT -3.750 747.800 -1.750 748.400 ;
        RECT -3.750 747.600 -1.950 747.800 ;
    END
  END WL703
  PIN WL704
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 746.150 -1.950 746.350 ;
        RECT -3.750 745.550 -1.750 746.150 ;
        RECT -3.750 745.350 -1.950 745.550 ;
    END
  END WL704
  PIN WL705
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 744.800 -1.950 745.000 ;
        RECT -3.750 744.200 -1.750 744.800 ;
        RECT -3.750 744.000 -1.950 744.200 ;
    END
  END WL705
  PIN WL706
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 742.550 -1.950 742.750 ;
        RECT -3.750 741.950 -1.750 742.550 ;
        RECT -3.750 741.750 -1.950 741.950 ;
    END
  END WL706
  PIN WL707
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 741.200 -1.950 741.400 ;
        RECT -3.750 740.600 -1.750 741.200 ;
        RECT -3.750 740.400 -1.950 740.600 ;
    END
  END WL707
  PIN WL708
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 738.950 -1.950 739.150 ;
        RECT -3.750 738.350 -1.750 738.950 ;
        RECT -3.750 738.150 -1.950 738.350 ;
    END
  END WL708
  PIN WL709
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 737.600 -1.950 737.800 ;
        RECT -3.750 737.000 -1.750 737.600 ;
        RECT -3.750 736.800 -1.950 737.000 ;
    END
  END WL709
  PIN WL710
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 735.350 -1.950 735.550 ;
        RECT -3.750 734.750 -1.750 735.350 ;
        RECT -3.750 734.550 -1.950 734.750 ;
    END
  END WL710
  PIN WL711
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 734.000 -1.950 734.200 ;
        RECT -3.750 733.400 -1.750 734.000 ;
        RECT -3.750 733.200 -1.950 733.400 ;
    END
  END WL711
  PIN WL712
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 731.750 -1.950 731.950 ;
        RECT -3.750 731.150 -1.750 731.750 ;
        RECT -3.750 730.950 -1.950 731.150 ;
    END
  END WL712
  PIN WL713
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 730.400 -1.950 730.600 ;
        RECT -3.750 729.800 -1.750 730.400 ;
        RECT -3.750 729.600 -1.950 729.800 ;
    END
  END WL713
  PIN WL714
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 728.150 -1.950 728.350 ;
        RECT -3.750 727.550 -1.750 728.150 ;
        RECT -3.750 727.350 -1.950 727.550 ;
    END
  END WL714
  PIN WL715
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 726.800 -1.950 727.000 ;
        RECT -3.750 726.200 -1.750 726.800 ;
        RECT -3.750 726.000 -1.950 726.200 ;
    END
  END WL715
  PIN WL716
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 724.550 -1.950 724.750 ;
        RECT -3.750 723.950 -1.750 724.550 ;
        RECT -3.750 723.750 -1.950 723.950 ;
    END
  END WL716
  PIN WL717
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 723.200 -1.950 723.400 ;
        RECT -3.750 722.600 -1.750 723.200 ;
        RECT -3.750 722.400 -1.950 722.600 ;
    END
  END WL717
  PIN WL718
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 720.950 -1.950 721.150 ;
        RECT -3.750 720.350 -1.750 720.950 ;
        RECT -3.750 720.150 -1.950 720.350 ;
    END
  END WL718
  PIN WL719
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 719.600 -1.950 719.800 ;
        RECT -3.750 719.000 -1.750 719.600 ;
        RECT -3.750 718.800 -1.950 719.000 ;
    END
  END WL719
  PIN WL720
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 717.350 -1.950 717.550 ;
        RECT -3.750 716.750 -1.750 717.350 ;
        RECT -3.750 716.550 -1.950 716.750 ;
    END
  END WL720
  PIN WL721
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 716.000 -1.950 716.200 ;
        RECT -3.750 715.400 -1.750 716.000 ;
        RECT -3.750 715.200 -1.950 715.400 ;
    END
  END WL721
  PIN WL722
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 713.750 -1.950 713.950 ;
        RECT -3.750 713.150 -1.750 713.750 ;
        RECT -3.750 712.950 -1.950 713.150 ;
    END
  END WL722
  PIN WL723
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 712.400 -1.950 712.600 ;
        RECT -3.750 711.800 -1.750 712.400 ;
        RECT -3.750 711.600 -1.950 711.800 ;
    END
  END WL723
  PIN WL724
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 710.150 -1.950 710.350 ;
        RECT -3.750 709.550 -1.750 710.150 ;
        RECT -3.750 709.350 -1.950 709.550 ;
    END
  END WL724
  PIN WL725
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 708.800 -1.950 709.000 ;
        RECT -3.750 708.200 -1.750 708.800 ;
        RECT -3.750 708.000 -1.950 708.200 ;
    END
  END WL725
  PIN WL726
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 706.550 -1.950 706.750 ;
        RECT -3.750 705.950 -1.750 706.550 ;
        RECT -3.750 705.750 -1.950 705.950 ;
    END
  END WL726
  PIN WL727
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 705.200 -1.950 705.400 ;
        RECT -3.750 704.600 -1.750 705.200 ;
        RECT -3.750 704.400 -1.950 704.600 ;
    END
  END WL727
  PIN WL728
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 702.950 -1.950 703.150 ;
        RECT -3.750 702.350 -1.750 702.950 ;
        RECT -3.750 702.150 -1.950 702.350 ;
    END
  END WL728
  PIN WL729
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 701.600 -1.950 701.800 ;
        RECT -3.750 701.000 -1.750 701.600 ;
        RECT -3.750 700.800 -1.950 701.000 ;
    END
  END WL729
  PIN WL730
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 699.350 -1.950 699.550 ;
        RECT -3.750 698.750 -1.750 699.350 ;
        RECT -3.750 698.550 -1.950 698.750 ;
    END
  END WL730
  PIN WL731
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 698.000 -1.950 698.200 ;
        RECT -3.750 697.400 -1.750 698.000 ;
        RECT -3.750 697.200 -1.950 697.400 ;
    END
  END WL731
  PIN WL732
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 695.750 -1.950 695.950 ;
        RECT -3.750 695.150 -1.750 695.750 ;
        RECT -3.750 694.950 -1.950 695.150 ;
    END
  END WL732
  PIN WL733
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 694.400 -1.950 694.600 ;
        RECT -3.750 693.800 -1.750 694.400 ;
        RECT -3.750 693.600 -1.950 693.800 ;
    END
  END WL733
  PIN WL734
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 692.150 -1.950 692.350 ;
        RECT -3.750 691.550 -1.750 692.150 ;
        RECT -3.750 691.350 -1.950 691.550 ;
    END
  END WL734
  PIN WL735
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 690.800 -1.950 691.000 ;
        RECT -3.750 690.200 -1.750 690.800 ;
        RECT -3.750 690.000 -1.950 690.200 ;
    END
  END WL735
  PIN WL736
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 688.550 -1.950 688.750 ;
        RECT -3.750 687.950 -1.750 688.550 ;
        RECT -3.750 687.750 -1.950 687.950 ;
    END
  END WL736
  PIN WL737
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 687.200 -1.950 687.400 ;
        RECT -3.750 686.600 -1.750 687.200 ;
        RECT -3.750 686.400 -1.950 686.600 ;
    END
  END WL737
  PIN WL738
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 684.950 -1.950 685.150 ;
        RECT -3.750 684.350 -1.750 684.950 ;
        RECT -3.750 684.150 -1.950 684.350 ;
    END
  END WL738
  PIN WL739
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 683.600 -1.950 683.800 ;
        RECT -3.750 683.000 -1.750 683.600 ;
        RECT -3.750 682.800 -1.950 683.000 ;
    END
  END WL739
  PIN WL740
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 681.350 -1.950 681.550 ;
        RECT -3.750 680.750 -1.750 681.350 ;
        RECT -3.750 680.550 -1.950 680.750 ;
    END
  END WL740
  PIN WL741
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 680.000 -1.950 680.200 ;
        RECT -3.750 679.400 -1.750 680.000 ;
        RECT -3.750 679.200 -1.950 679.400 ;
    END
  END WL741
  PIN WL742
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 677.750 -1.950 677.950 ;
        RECT -3.750 677.150 -1.750 677.750 ;
        RECT -3.750 676.950 -1.950 677.150 ;
    END
  END WL742
  PIN WL743
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 676.400 -1.950 676.600 ;
        RECT -3.750 675.800 -1.750 676.400 ;
        RECT -3.750 675.600 -1.950 675.800 ;
    END
  END WL743
  PIN WL744
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 674.150 -1.950 674.350 ;
        RECT -3.750 673.550 -1.750 674.150 ;
        RECT -3.750 673.350 -1.950 673.550 ;
    END
  END WL744
  PIN WL745
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 672.800 -1.950 673.000 ;
        RECT -3.750 672.200 -1.750 672.800 ;
        RECT -3.750 672.000 -1.950 672.200 ;
    END
  END WL745
  PIN WL746
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 670.550 -1.950 670.750 ;
        RECT -3.750 669.950 -1.750 670.550 ;
        RECT -3.750 669.750 -1.950 669.950 ;
    END
  END WL746
  PIN WL747
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 669.200 -1.950 669.400 ;
        RECT -3.750 668.600 -1.750 669.200 ;
        RECT -3.750 668.400 -1.950 668.600 ;
    END
  END WL747
  PIN WL748
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 666.950 -1.950 667.150 ;
        RECT -3.750 666.350 -1.750 666.950 ;
        RECT -3.750 666.150 -1.950 666.350 ;
    END
  END WL748
  PIN WL749
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 665.600 -1.950 665.800 ;
        RECT -3.750 665.000 -1.750 665.600 ;
        RECT -3.750 664.800 -1.950 665.000 ;
    END
  END WL749
  PIN WL750
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 663.350 -1.950 663.550 ;
        RECT -3.750 662.750 -1.750 663.350 ;
        RECT -3.750 662.550 -1.950 662.750 ;
    END
  END WL750
  PIN WL751
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 662.000 -1.950 662.200 ;
        RECT -3.750 661.400 -1.750 662.000 ;
        RECT -3.750 661.200 -1.950 661.400 ;
    END
  END WL751
  PIN WL752
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 659.750 -1.950 659.950 ;
        RECT -3.750 659.150 -1.750 659.750 ;
        RECT -3.750 658.950 -1.950 659.150 ;
    END
  END WL752
  PIN WL753
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 658.400 -1.950 658.600 ;
        RECT -3.750 657.800 -1.750 658.400 ;
        RECT -3.750 657.600 -1.950 657.800 ;
    END
  END WL753
  PIN WL754
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 656.150 -1.950 656.350 ;
        RECT -3.750 655.550 -1.750 656.150 ;
        RECT -3.750 655.350 -1.950 655.550 ;
    END
  END WL754
  PIN WL755
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 654.800 -1.950 655.000 ;
        RECT -3.750 654.200 -1.750 654.800 ;
        RECT -3.750 654.000 -1.950 654.200 ;
    END
  END WL755
  PIN WL756
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 652.550 -1.950 652.750 ;
        RECT -3.750 651.950 -1.750 652.550 ;
        RECT -3.750 651.750 -1.950 651.950 ;
    END
  END WL756
  PIN WL757
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 651.200 -1.950 651.400 ;
        RECT -3.750 650.600 -1.750 651.200 ;
        RECT -3.750 650.400 -1.950 650.600 ;
    END
  END WL757
  PIN WL758
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 648.950 -1.950 649.150 ;
        RECT -3.750 648.350 -1.750 648.950 ;
        RECT -3.750 648.150 -1.950 648.350 ;
    END
  END WL758
  PIN WL759
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 647.600 -1.950 647.800 ;
        RECT -3.750 647.000 -1.750 647.600 ;
        RECT -3.750 646.800 -1.950 647.000 ;
    END
  END WL759
  PIN WL760
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 645.350 -1.950 645.550 ;
        RECT -3.750 644.750 -1.750 645.350 ;
        RECT -3.750 644.550 -1.950 644.750 ;
    END
  END WL760
  PIN WL761
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 644.000 -1.950 644.200 ;
        RECT -3.750 643.400 -1.750 644.000 ;
        RECT -3.750 643.200 -1.950 643.400 ;
    END
  END WL761
  PIN WL762
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 641.750 -1.950 641.950 ;
        RECT -3.750 641.150 -1.750 641.750 ;
        RECT -3.750 640.950 -1.950 641.150 ;
    END
  END WL762
  PIN WL763
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 640.400 -1.950 640.600 ;
        RECT -3.750 639.800 -1.750 640.400 ;
        RECT -3.750 639.600 -1.950 639.800 ;
    END
  END WL763
  PIN WL764
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 638.150 -1.950 638.350 ;
        RECT -3.750 637.550 -1.750 638.150 ;
        RECT -3.750 637.350 -1.950 637.550 ;
    END
  END WL764
  PIN WL765
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 636.800 -1.950 637.000 ;
        RECT -3.750 636.200 -1.750 636.800 ;
        RECT -3.750 636.000 -1.950 636.200 ;
    END
  END WL765
  PIN WL766
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 634.550 -1.950 634.750 ;
        RECT -3.750 633.950 -1.750 634.550 ;
        RECT -3.750 633.750 -1.950 633.950 ;
    END
  END WL766
  PIN WL767
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 633.200 -1.950 633.400 ;
        RECT -3.750 632.600 -1.750 633.200 ;
        RECT -3.750 632.400 -1.950 632.600 ;
    END
  END WL767
  PIN WL768
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 630.950 -1.950 631.150 ;
        RECT -3.750 630.350 -1.750 630.950 ;
        RECT -3.750 630.150 -1.950 630.350 ;
    END
  END WL768
  PIN WL769
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 629.600 -1.950 629.800 ;
        RECT -3.750 629.000 -1.750 629.600 ;
        RECT -3.750 628.800 -1.950 629.000 ;
    END
  END WL769
  PIN WL770
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 627.350 -1.950 627.550 ;
        RECT -3.750 626.750 -1.750 627.350 ;
        RECT -3.750 626.550 -1.950 626.750 ;
    END
  END WL770
  PIN WL771
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 626.000 -1.950 626.200 ;
        RECT -3.750 625.400 -1.750 626.000 ;
        RECT -3.750 625.200 -1.950 625.400 ;
    END
  END WL771
  PIN WL772
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 623.750 -1.950 623.950 ;
        RECT -3.750 623.150 -1.750 623.750 ;
        RECT -3.750 622.950 -1.950 623.150 ;
    END
  END WL772
  PIN WL773
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 622.400 -1.950 622.600 ;
        RECT -3.750 621.800 -1.750 622.400 ;
        RECT -3.750 621.600 -1.950 621.800 ;
    END
  END WL773
  PIN WL774
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 619.600 -1.950 619.800 ;
        RECT -3.750 619.000 -1.750 619.600 ;
        RECT -3.750 618.800 -1.950 619.000 ;
    END
  END WL774
  PIN WL775
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 618.250 -1.950 618.450 ;
        RECT -3.750 617.650 -1.750 618.250 ;
        RECT -3.750 617.450 -1.950 617.650 ;
    END
  END WL775
  PIN WL776
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 616.000 -1.950 616.200 ;
        RECT -3.750 615.400 -1.750 616.000 ;
        RECT -3.750 615.200 -1.950 615.400 ;
    END
  END WL776
  PIN WL777
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 614.650 -1.950 614.850 ;
        RECT -3.750 614.050 -1.750 614.650 ;
        RECT -3.750 613.850 -1.950 614.050 ;
    END
  END WL777
  PIN WL778
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 612.400 -1.950 612.600 ;
        RECT -3.750 611.800 -1.750 612.400 ;
        RECT -3.750 611.600 -1.950 611.800 ;
    END
  END WL778
  PIN WL779
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 611.050 -1.950 611.250 ;
        RECT -3.750 610.450 -1.750 611.050 ;
        RECT -3.750 610.250 -1.950 610.450 ;
    END
  END WL779
  PIN WL780
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 608.800 -1.950 609.000 ;
        RECT -3.750 608.200 -1.750 608.800 ;
        RECT -3.750 608.000 -1.950 608.200 ;
    END
  END WL780
  PIN WL781
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 607.450 -1.950 607.650 ;
        RECT -3.750 606.850 -1.750 607.450 ;
        RECT -3.750 606.650 -1.950 606.850 ;
    END
  END WL781
  PIN WL782
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 605.200 -1.950 605.400 ;
        RECT -3.750 604.600 -1.750 605.200 ;
        RECT -3.750 604.400 -1.950 604.600 ;
    END
  END WL782
  PIN WL783
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 603.850 -1.950 604.050 ;
        RECT -3.750 603.250 -1.750 603.850 ;
        RECT -3.750 603.050 -1.950 603.250 ;
    END
  END WL783
  PIN WL784
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 601.600 -1.950 601.800 ;
        RECT -3.750 601.000 -1.750 601.600 ;
        RECT -3.750 600.800 -1.950 601.000 ;
    END
  END WL784
  PIN WL785
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 600.250 -1.950 600.450 ;
        RECT -3.750 599.650 -1.750 600.250 ;
        RECT -3.750 599.450 -1.950 599.650 ;
    END
  END WL785
  PIN WL786
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 598.000 -1.950 598.200 ;
        RECT -3.750 597.400 -1.750 598.000 ;
        RECT -3.750 597.200 -1.950 597.400 ;
    END
  END WL786
  PIN WL787
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 596.650 -1.950 596.850 ;
        RECT -3.750 596.050 -1.750 596.650 ;
        RECT -3.750 595.850 -1.950 596.050 ;
    END
  END WL787
  PIN WL788
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 594.400 -1.950 594.600 ;
        RECT -3.750 593.800 -1.750 594.400 ;
        RECT -3.750 593.600 -1.950 593.800 ;
    END
  END WL788
  PIN WL789
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 593.050 -1.950 593.250 ;
        RECT -3.750 592.450 -1.750 593.050 ;
        RECT -3.750 592.250 -1.950 592.450 ;
    END
  END WL789
  PIN WL790
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 590.800 -1.950 591.000 ;
        RECT -3.750 590.200 -1.750 590.800 ;
        RECT -3.750 590.000 -1.950 590.200 ;
    END
  END WL790
  PIN WL791
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 589.450 -1.950 589.650 ;
        RECT -3.750 588.850 -1.750 589.450 ;
        RECT -3.750 588.650 -1.950 588.850 ;
    END
  END WL791
  PIN WL792
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 587.200 -1.950 587.400 ;
        RECT -3.750 586.600 -1.750 587.200 ;
        RECT -3.750 586.400 -1.950 586.600 ;
    END
  END WL792
  PIN WL793
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 585.850 -1.950 586.050 ;
        RECT -3.750 585.250 -1.750 585.850 ;
        RECT -3.750 585.050 -1.950 585.250 ;
    END
  END WL793
  PIN WL794
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 583.600 -1.950 583.800 ;
        RECT -3.750 583.000 -1.750 583.600 ;
        RECT -3.750 582.800 -1.950 583.000 ;
    END
  END WL794
  PIN WL795
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 582.250 -1.950 582.450 ;
        RECT -3.750 581.650 -1.750 582.250 ;
        RECT -3.750 581.450 -1.950 581.650 ;
    END
  END WL795
  PIN WL796
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 580.000 -1.950 580.200 ;
        RECT -3.750 579.400 -1.750 580.000 ;
        RECT -3.750 579.200 -1.950 579.400 ;
    END
  END WL796
  PIN WL797
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 578.650 -1.950 578.850 ;
        RECT -3.750 578.050 -1.750 578.650 ;
        RECT -3.750 577.850 -1.950 578.050 ;
    END
  END WL797
  PIN WL798
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 576.400 -1.950 576.600 ;
        RECT -3.750 575.800 -1.750 576.400 ;
        RECT -3.750 575.600 -1.950 575.800 ;
    END
  END WL798
  PIN WL799
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 575.050 -1.950 575.250 ;
        RECT -3.750 574.450 -1.750 575.050 ;
        RECT -3.750 574.250 -1.950 574.450 ;
    END
  END WL799
  PIN WL800
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 572.800 -1.950 573.000 ;
        RECT -3.750 572.200 -1.750 572.800 ;
        RECT -3.750 572.000 -1.950 572.200 ;
    END
  END WL800
  PIN WL801
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 571.450 -1.950 571.650 ;
        RECT -3.750 570.850 -1.750 571.450 ;
        RECT -3.750 570.650 -1.950 570.850 ;
    END
  END WL801
  PIN WL802
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 569.200 -1.950 569.400 ;
        RECT -3.750 568.600 -1.750 569.200 ;
        RECT -3.750 568.400 -1.950 568.600 ;
    END
  END WL802
  PIN WL803
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 567.850 -1.950 568.050 ;
        RECT -3.750 567.250 -1.750 567.850 ;
        RECT -3.750 567.050 -1.950 567.250 ;
    END
  END WL803
  PIN WL804
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 565.600 -1.950 565.800 ;
        RECT -3.750 565.000 -1.750 565.600 ;
        RECT -3.750 564.800 -1.950 565.000 ;
    END
  END WL804
  PIN WL805
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 564.250 -1.950 564.450 ;
        RECT -3.750 563.650 -1.750 564.250 ;
        RECT -3.750 563.450 -1.950 563.650 ;
    END
  END WL805
  PIN WL806
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 562.000 -1.950 562.200 ;
        RECT -3.750 561.400 -1.750 562.000 ;
        RECT -3.750 561.200 -1.950 561.400 ;
    END
  END WL806
  PIN WL807
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 560.650 -1.950 560.850 ;
        RECT -3.750 560.050 -1.750 560.650 ;
        RECT -3.750 559.850 -1.950 560.050 ;
    END
  END WL807
  PIN WL808
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 558.400 -1.950 558.600 ;
        RECT -3.750 557.800 -1.750 558.400 ;
        RECT -3.750 557.600 -1.950 557.800 ;
    END
  END WL808
  PIN WL809
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 557.050 -1.950 557.250 ;
        RECT -3.750 556.450 -1.750 557.050 ;
        RECT -3.750 556.250 -1.950 556.450 ;
    END
  END WL809
  PIN WL810
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 554.800 -1.950 555.000 ;
        RECT -3.750 554.200 -1.750 554.800 ;
        RECT -3.750 554.000 -1.950 554.200 ;
    END
  END WL810
  PIN WL811
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 553.450 -1.950 553.650 ;
        RECT -3.750 552.850 -1.750 553.450 ;
        RECT -3.750 552.650 -1.950 552.850 ;
    END
  END WL811
  PIN WL812
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 551.200 -1.950 551.400 ;
        RECT -3.750 550.600 -1.750 551.200 ;
        RECT -3.750 550.400 -1.950 550.600 ;
    END
  END WL812
  PIN WL813
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 549.850 -1.950 550.050 ;
        RECT -3.750 549.250 -1.750 549.850 ;
        RECT -3.750 549.050 -1.950 549.250 ;
    END
  END WL813
  PIN WL814
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 547.600 -1.950 547.800 ;
        RECT -3.750 547.000 -1.750 547.600 ;
        RECT -3.750 546.800 -1.950 547.000 ;
    END
  END WL814
  PIN WL815
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 546.250 -1.950 546.450 ;
        RECT -3.750 545.650 -1.750 546.250 ;
        RECT -3.750 545.450 -1.950 545.650 ;
    END
  END WL815
  PIN WL816
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 544.000 -1.950 544.200 ;
        RECT -3.750 543.400 -1.750 544.000 ;
        RECT -3.750 543.200 -1.950 543.400 ;
    END
  END WL816
  PIN WL817
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 542.650 -1.950 542.850 ;
        RECT -3.750 542.050 -1.750 542.650 ;
        RECT -3.750 541.850 -1.950 542.050 ;
    END
  END WL817
  PIN WL818
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 540.400 -1.950 540.600 ;
        RECT -3.750 539.800 -1.750 540.400 ;
        RECT -3.750 539.600 -1.950 539.800 ;
    END
  END WL818
  PIN WL819
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 539.050 -1.950 539.250 ;
        RECT -3.750 538.450 -1.750 539.050 ;
        RECT -3.750 538.250 -1.950 538.450 ;
    END
  END WL819
  PIN WL820
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 536.800 -1.950 537.000 ;
        RECT -3.750 536.200 -1.750 536.800 ;
        RECT -3.750 536.000 -1.950 536.200 ;
    END
  END WL820
  PIN WL821
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 535.450 -1.950 535.650 ;
        RECT -3.750 534.850 -1.750 535.450 ;
        RECT -3.750 534.650 -1.950 534.850 ;
    END
  END WL821
  PIN WL822
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 533.200 -1.950 533.400 ;
        RECT -3.750 532.600 -1.750 533.200 ;
        RECT -3.750 532.400 -1.950 532.600 ;
    END
  END WL822
  PIN WL823
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 531.850 -1.950 532.050 ;
        RECT -3.750 531.250 -1.750 531.850 ;
        RECT -3.750 531.050 -1.950 531.250 ;
    END
  END WL823
  PIN WL824
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 529.600 -1.950 529.800 ;
        RECT -3.750 529.000 -1.750 529.600 ;
        RECT -3.750 528.800 -1.950 529.000 ;
    END
  END WL824
  PIN WL825
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 528.250 -1.950 528.450 ;
        RECT -3.750 527.650 -1.750 528.250 ;
        RECT -3.750 527.450 -1.950 527.650 ;
    END
  END WL825
  PIN WL826
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 526.000 -1.950 526.200 ;
        RECT -3.750 525.400 -1.750 526.000 ;
        RECT -3.750 525.200 -1.950 525.400 ;
    END
  END WL826
  PIN WL827
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 524.650 -1.950 524.850 ;
        RECT -3.750 524.050 -1.750 524.650 ;
        RECT -3.750 523.850 -1.950 524.050 ;
    END
  END WL827
  PIN WL828
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 522.400 -1.950 522.600 ;
        RECT -3.750 521.800 -1.750 522.400 ;
        RECT -3.750 521.600 -1.950 521.800 ;
    END
  END WL828
  PIN WL829
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 521.050 -1.950 521.250 ;
        RECT -3.750 520.450 -1.750 521.050 ;
        RECT -3.750 520.250 -1.950 520.450 ;
    END
  END WL829
  PIN WL830
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 518.800 -1.950 519.000 ;
        RECT -3.750 518.200 -1.750 518.800 ;
        RECT -3.750 518.000 -1.950 518.200 ;
    END
  END WL830
  PIN WL831
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 517.450 -1.950 517.650 ;
        RECT -3.750 516.850 -1.750 517.450 ;
        RECT -3.750 516.650 -1.950 516.850 ;
    END
  END WL831
  PIN WL832
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 515.200 -1.950 515.400 ;
        RECT -3.750 514.600 -1.750 515.200 ;
        RECT -3.750 514.400 -1.950 514.600 ;
    END
  END WL832
  PIN WL833
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 513.850 -1.950 514.050 ;
        RECT -3.750 513.250 -1.750 513.850 ;
        RECT -3.750 513.050 -1.950 513.250 ;
    END
  END WL833
  PIN WL834
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 511.600 -1.950 511.800 ;
        RECT -3.750 511.000 -1.750 511.600 ;
        RECT -3.750 510.800 -1.950 511.000 ;
    END
  END WL834
  PIN WL835
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 510.250 -1.950 510.450 ;
        RECT -3.750 509.650 -1.750 510.250 ;
        RECT -3.750 509.450 -1.950 509.650 ;
    END
  END WL835
  PIN WL836
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 508.000 -1.950 508.200 ;
        RECT -3.750 507.400 -1.750 508.000 ;
        RECT -3.750 507.200 -1.950 507.400 ;
    END
  END WL836
  PIN WL837
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 506.650 -1.950 506.850 ;
        RECT -3.750 506.050 -1.750 506.650 ;
        RECT -3.750 505.850 -1.950 506.050 ;
    END
  END WL837
  PIN WL838
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 504.400 -1.950 504.600 ;
        RECT -3.750 503.800 -1.750 504.400 ;
        RECT -3.750 503.600 -1.950 503.800 ;
    END
  END WL838
  PIN WL839
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 503.050 -1.950 503.250 ;
        RECT -3.750 502.450 -1.750 503.050 ;
        RECT -3.750 502.250 -1.950 502.450 ;
    END
  END WL839
  PIN WL840
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 500.800 -1.950 501.000 ;
        RECT -3.750 500.200 -1.750 500.800 ;
        RECT -3.750 500.000 -1.950 500.200 ;
    END
  END WL840
  PIN WL841
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 499.450 -1.950 499.650 ;
        RECT -3.750 498.850 -1.750 499.450 ;
        RECT -3.750 498.650 -1.950 498.850 ;
    END
  END WL841
  PIN WL842
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 497.200 -1.950 497.400 ;
        RECT -3.750 496.600 -1.750 497.200 ;
        RECT -3.750 496.400 -1.950 496.600 ;
    END
  END WL842
  PIN WL843
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 495.850 -1.950 496.050 ;
        RECT -3.750 495.250 -1.750 495.850 ;
        RECT -3.750 495.050 -1.950 495.250 ;
    END
  END WL843
  PIN WL844
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 493.600 -1.950 493.800 ;
        RECT -3.750 493.000 -1.750 493.600 ;
        RECT -3.750 492.800 -1.950 493.000 ;
    END
  END WL844
  PIN WL845
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 492.250 -1.950 492.450 ;
        RECT -3.750 491.650 -1.750 492.250 ;
        RECT -3.750 491.450 -1.950 491.650 ;
    END
  END WL845
  PIN WL846
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 490.000 -1.950 490.200 ;
        RECT -3.750 489.400 -1.750 490.000 ;
        RECT -3.750 489.200 -1.950 489.400 ;
    END
  END WL846
  PIN WL847
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 488.650 -1.950 488.850 ;
        RECT -3.750 488.050 -1.750 488.650 ;
        RECT -3.750 487.850 -1.950 488.050 ;
    END
  END WL847
  PIN WL848
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 486.400 -1.950 486.600 ;
        RECT -3.750 485.800 -1.750 486.400 ;
        RECT -3.750 485.600 -1.950 485.800 ;
    END
  END WL848
  PIN WL849
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 485.050 -1.950 485.250 ;
        RECT -3.750 484.450 -1.750 485.050 ;
        RECT -3.750 484.250 -1.950 484.450 ;
    END
  END WL849
  PIN WL850
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 482.800 -1.950 483.000 ;
        RECT -3.750 482.200 -1.750 482.800 ;
        RECT -3.750 482.000 -1.950 482.200 ;
    END
  END WL850
  PIN WL851
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 481.450 -1.950 481.650 ;
        RECT -3.750 480.850 -1.750 481.450 ;
        RECT -3.750 480.650 -1.950 480.850 ;
    END
  END WL851
  PIN WL852
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 479.200 -1.950 479.400 ;
        RECT -3.750 478.600 -1.750 479.200 ;
        RECT -3.750 478.400 -1.950 478.600 ;
    END
  END WL852
  PIN WL853
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 477.850 -1.950 478.050 ;
        RECT -3.750 477.250 -1.750 477.850 ;
        RECT -3.750 477.050 -1.950 477.250 ;
    END
  END WL853
  PIN WL854
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 475.600 -1.950 475.800 ;
        RECT -3.750 475.000 -1.750 475.600 ;
        RECT -3.750 474.800 -1.950 475.000 ;
    END
  END WL854
  PIN WL855
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 474.250 -1.950 474.450 ;
        RECT -3.750 473.650 -1.750 474.250 ;
        RECT -3.750 473.450 -1.950 473.650 ;
    END
  END WL855
  PIN WL856
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 472.000 -1.950 472.200 ;
        RECT -3.750 471.400 -1.750 472.000 ;
        RECT -3.750 471.200 -1.950 471.400 ;
    END
  END WL856
  PIN WL857
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 470.650 -1.950 470.850 ;
        RECT -3.750 470.050 -1.750 470.650 ;
        RECT -3.750 469.850 -1.950 470.050 ;
    END
  END WL857
  PIN WL858
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 468.400 -1.950 468.600 ;
        RECT -3.750 467.800 -1.750 468.400 ;
        RECT -3.750 467.600 -1.950 467.800 ;
    END
  END WL858
  PIN WL859
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 467.050 -1.950 467.250 ;
        RECT -3.750 466.450 -1.750 467.050 ;
        RECT -3.750 466.250 -1.950 466.450 ;
    END
  END WL859
  PIN WL860
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 464.800 -1.950 465.000 ;
        RECT -3.750 464.200 -1.750 464.800 ;
        RECT -3.750 464.000 -1.950 464.200 ;
    END
  END WL860
  PIN WL861
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 463.450 -1.950 463.650 ;
        RECT -3.750 462.850 -1.750 463.450 ;
        RECT -3.750 462.650 -1.950 462.850 ;
    END
  END WL861
  PIN WL862
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 461.200 -1.950 461.400 ;
        RECT -3.750 460.600 -1.750 461.200 ;
        RECT -3.750 460.400 -1.950 460.600 ;
    END
  END WL862
  PIN WL863
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 459.850 -1.950 460.050 ;
        RECT -3.750 459.250 -1.750 459.850 ;
        RECT -3.750 459.050 -1.950 459.250 ;
    END
  END WL863
  PIN WL864
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 457.600 -1.950 457.800 ;
        RECT -3.750 457.000 -1.750 457.600 ;
        RECT -3.750 456.800 -1.950 457.000 ;
    END
  END WL864
  PIN WL865
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 456.250 -1.950 456.450 ;
        RECT -3.750 455.650 -1.750 456.250 ;
        RECT -3.750 455.450 -1.950 455.650 ;
    END
  END WL865
  PIN WL866
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 454.000 -1.950 454.200 ;
        RECT -3.750 453.400 -1.750 454.000 ;
        RECT -3.750 453.200 -1.950 453.400 ;
    END
  END WL866
  PIN WL867
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 452.650 -1.950 452.850 ;
        RECT -3.750 452.050 -1.750 452.650 ;
        RECT -3.750 451.850 -1.950 452.050 ;
    END
  END WL867
  PIN WL868
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 450.400 -1.950 450.600 ;
        RECT -3.750 449.800 -1.750 450.400 ;
        RECT -3.750 449.600 -1.950 449.800 ;
    END
  END WL868
  PIN WL869
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 449.050 -1.950 449.250 ;
        RECT -3.750 448.450 -1.750 449.050 ;
        RECT -3.750 448.250 -1.950 448.450 ;
    END
  END WL869
  PIN WL870
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 446.800 -1.950 447.000 ;
        RECT -3.750 446.200 -1.750 446.800 ;
        RECT -3.750 446.000 -1.950 446.200 ;
    END
  END WL870
  PIN WL871
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 445.450 -1.950 445.650 ;
        RECT -3.750 444.850 -1.750 445.450 ;
        RECT -3.750 444.650 -1.950 444.850 ;
    END
  END WL871
  PIN WL872
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 443.200 -1.950 443.400 ;
        RECT -3.750 442.600 -1.750 443.200 ;
        RECT -3.750 442.400 -1.950 442.600 ;
    END
  END WL872
  PIN WL873
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 441.850 -1.950 442.050 ;
        RECT -3.750 441.250 -1.750 441.850 ;
        RECT -3.750 441.050 -1.950 441.250 ;
    END
  END WL873
  PIN WL874
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 439.600 -1.950 439.800 ;
        RECT -3.750 439.000 -1.750 439.600 ;
        RECT -3.750 438.800 -1.950 439.000 ;
    END
  END WL874
  PIN WL875
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 438.250 -1.950 438.450 ;
        RECT -3.750 437.650 -1.750 438.250 ;
        RECT -3.750 437.450 -1.950 437.650 ;
    END
  END WL875
  PIN WL876
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 436.000 -1.950 436.200 ;
        RECT -3.750 435.400 -1.750 436.000 ;
        RECT -3.750 435.200 -1.950 435.400 ;
    END
  END WL876
  PIN WL877
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 434.650 -1.950 434.850 ;
        RECT -3.750 434.050 -1.750 434.650 ;
        RECT -3.750 433.850 -1.950 434.050 ;
    END
  END WL877
  PIN WL878
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 432.400 -1.950 432.600 ;
        RECT -3.750 431.800 -1.750 432.400 ;
        RECT -3.750 431.600 -1.950 431.800 ;
    END
  END WL878
  PIN WL879
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 431.050 -1.950 431.250 ;
        RECT -3.750 430.450 -1.750 431.050 ;
        RECT -3.750 430.250 -1.950 430.450 ;
    END
  END WL879
  PIN WL880
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 428.800 -1.950 429.000 ;
        RECT -3.750 428.200 -1.750 428.800 ;
        RECT -3.750 428.000 -1.950 428.200 ;
    END
  END WL880
  PIN WL881
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 427.450 -1.950 427.650 ;
        RECT -3.750 426.850 -1.750 427.450 ;
        RECT -3.750 426.650 -1.950 426.850 ;
    END
  END WL881
  PIN WL882
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 425.200 -1.950 425.400 ;
        RECT -3.750 424.600 -1.750 425.200 ;
        RECT -3.750 424.400 -1.950 424.600 ;
    END
  END WL882
  PIN WL883
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 423.850 -1.950 424.050 ;
        RECT -3.750 423.250 -1.750 423.850 ;
        RECT -3.750 423.050 -1.950 423.250 ;
    END
  END WL883
  PIN WL884
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 421.050 -1.950 421.250 ;
        RECT -3.750 420.450 -1.750 421.050 ;
        RECT -3.750 420.250 -1.950 420.450 ;
    END
  END WL884
  PIN WL885
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 419.700 -1.950 419.900 ;
        RECT -3.750 419.100 -1.750 419.700 ;
        RECT -3.750 418.900 -1.950 419.100 ;
    END
  END WL885
  PIN WL886
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 417.450 -1.950 417.650 ;
        RECT -3.750 416.850 -1.750 417.450 ;
        RECT -3.750 416.650 -1.950 416.850 ;
    END
  END WL886
  PIN WL887
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 416.100 -1.950 416.300 ;
        RECT -3.750 415.500 -1.750 416.100 ;
        RECT -3.750 415.300 -1.950 415.500 ;
    END
  END WL887
  PIN WL888
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 413.850 -1.950 414.050 ;
        RECT -3.750 413.250 -1.750 413.850 ;
        RECT -3.750 413.050 -1.950 413.250 ;
    END
  END WL888
  PIN WL889
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 412.500 -1.950 412.700 ;
        RECT -3.750 411.900 -1.750 412.500 ;
        RECT -3.750 411.700 -1.950 411.900 ;
    END
  END WL889
  PIN WL890
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 410.250 -1.950 410.450 ;
        RECT -3.750 409.650 -1.750 410.250 ;
        RECT -3.750 409.450 -1.950 409.650 ;
    END
  END WL890
  PIN WL891
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 408.900 -1.950 409.100 ;
        RECT -3.750 408.300 -1.750 408.900 ;
        RECT -3.750 408.100 -1.950 408.300 ;
    END
  END WL891
  PIN WL892
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 406.650 -1.950 406.850 ;
        RECT -3.750 406.050 -1.750 406.650 ;
        RECT -3.750 405.850 -1.950 406.050 ;
    END
  END WL892
  PIN WL893
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 405.300 -1.950 405.500 ;
        RECT -3.750 404.700 -1.750 405.300 ;
        RECT -3.750 404.500 -1.950 404.700 ;
    END
  END WL893
  PIN WL894
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 403.050 -1.950 403.250 ;
        RECT -3.750 402.450 -1.750 403.050 ;
        RECT -3.750 402.250 -1.950 402.450 ;
    END
  END WL894
  PIN WL895
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 401.700 -1.950 401.900 ;
        RECT -3.750 401.100 -1.750 401.700 ;
        RECT -3.750 400.900 -1.950 401.100 ;
    END
  END WL895
  PIN WL896
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 399.450 -1.950 399.650 ;
        RECT -3.750 398.850 -1.750 399.450 ;
        RECT -3.750 398.650 -1.950 398.850 ;
    END
  END WL896
  PIN WL897
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 398.100 -1.950 398.300 ;
        RECT -3.750 397.500 -1.750 398.100 ;
        RECT -3.750 397.300 -1.950 397.500 ;
    END
  END WL897
  PIN WL898
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 395.850 -1.950 396.050 ;
        RECT -3.750 395.250 -1.750 395.850 ;
        RECT -3.750 395.050 -1.950 395.250 ;
    END
  END WL898
  PIN WL899
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 394.500 -1.950 394.700 ;
        RECT -3.750 393.900 -1.750 394.500 ;
        RECT -3.750 393.700 -1.950 393.900 ;
    END
  END WL899
  PIN WL900
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 392.250 -1.950 392.450 ;
        RECT -3.750 391.650 -1.750 392.250 ;
        RECT -3.750 391.450 -1.950 391.650 ;
    END
  END WL900
  PIN WL901
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 390.900 -1.950 391.100 ;
        RECT -3.750 390.300 -1.750 390.900 ;
        RECT -3.750 390.100 -1.950 390.300 ;
    END
  END WL901
  PIN WL902
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 388.650 -1.950 388.850 ;
        RECT -3.750 388.050 -1.750 388.650 ;
        RECT -3.750 387.850 -1.950 388.050 ;
    END
  END WL902
  PIN WL903
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 387.300 -1.950 387.500 ;
        RECT -3.750 386.700 -1.750 387.300 ;
        RECT -3.750 386.500 -1.950 386.700 ;
    END
  END WL903
  PIN WL904
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 385.050 -1.950 385.250 ;
        RECT -3.750 384.450 -1.750 385.050 ;
        RECT -3.750 384.250 -1.950 384.450 ;
    END
  END WL904
  PIN WL905
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 383.700 -1.950 383.900 ;
        RECT -3.750 383.100 -1.750 383.700 ;
        RECT -3.750 382.900 -1.950 383.100 ;
    END
  END WL905
  PIN WL906
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 381.450 -1.950 381.650 ;
        RECT -3.750 380.850 -1.750 381.450 ;
        RECT -3.750 380.650 -1.950 380.850 ;
    END
  END WL906
  PIN WL907
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 380.100 -1.950 380.300 ;
        RECT -3.750 379.500 -1.750 380.100 ;
        RECT -3.750 379.300 -1.950 379.500 ;
    END
  END WL907
  PIN WL908
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 377.850 -1.950 378.050 ;
        RECT -3.750 377.250 -1.750 377.850 ;
        RECT -3.750 377.050 -1.950 377.250 ;
    END
  END WL908
  PIN WL909
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 376.500 -1.950 376.700 ;
        RECT -3.750 375.900 -1.750 376.500 ;
        RECT -3.750 375.700 -1.950 375.900 ;
    END
  END WL909
  PIN WL910
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 374.250 -1.950 374.450 ;
        RECT -3.750 373.650 -1.750 374.250 ;
        RECT -3.750 373.450 -1.950 373.650 ;
    END
  END WL910
  PIN WL911
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 372.900 -1.950 373.100 ;
        RECT -3.750 372.300 -1.750 372.900 ;
        RECT -3.750 372.100 -1.950 372.300 ;
    END
  END WL911
  PIN WL912
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 370.650 -1.950 370.850 ;
        RECT -3.750 370.050 -1.750 370.650 ;
        RECT -3.750 369.850 -1.950 370.050 ;
    END
  END WL912
  PIN WL913
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 369.300 -1.950 369.500 ;
        RECT -3.750 368.700 -1.750 369.300 ;
        RECT -3.750 368.500 -1.950 368.700 ;
    END
  END WL913
  PIN WL914
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 367.050 -1.950 367.250 ;
        RECT -3.750 366.450 -1.750 367.050 ;
        RECT -3.750 366.250 -1.950 366.450 ;
    END
  END WL914
  PIN WL915
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 365.700 -1.950 365.900 ;
        RECT -3.750 365.100 -1.750 365.700 ;
        RECT -3.750 364.900 -1.950 365.100 ;
    END
  END WL915
  PIN WL916
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 363.450 -1.950 363.650 ;
        RECT -3.750 362.850 -1.750 363.450 ;
        RECT -3.750 362.650 -1.950 362.850 ;
    END
  END WL916
  PIN WL917
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 362.100 -1.950 362.300 ;
        RECT -3.750 361.500 -1.750 362.100 ;
        RECT -3.750 361.300 -1.950 361.500 ;
    END
  END WL917
  PIN WL918
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 359.850 -1.950 360.050 ;
        RECT -3.750 359.250 -1.750 359.850 ;
        RECT -3.750 359.050 -1.950 359.250 ;
    END
  END WL918
  PIN WL919
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 358.500 -1.950 358.700 ;
        RECT -3.750 357.900 -1.750 358.500 ;
        RECT -3.750 357.700 -1.950 357.900 ;
    END
  END WL919
  PIN WL920
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 356.250 -1.950 356.450 ;
        RECT -3.750 355.650 -1.750 356.250 ;
        RECT -3.750 355.450 -1.950 355.650 ;
    END
  END WL920
  PIN WL921
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 354.900 -1.950 355.100 ;
        RECT -3.750 354.300 -1.750 354.900 ;
        RECT -3.750 354.100 -1.950 354.300 ;
    END
  END WL921
  PIN WL922
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 352.650 -1.950 352.850 ;
        RECT -3.750 352.050 -1.750 352.650 ;
        RECT -3.750 351.850 -1.950 352.050 ;
    END
  END WL922
  PIN WL923
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 351.300 -1.950 351.500 ;
        RECT -3.750 350.700 -1.750 351.300 ;
        RECT -3.750 350.500 -1.950 350.700 ;
    END
  END WL923
  PIN WL924
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 349.050 -1.950 349.250 ;
        RECT -3.750 348.450 -1.750 349.050 ;
        RECT -3.750 348.250 -1.950 348.450 ;
    END
  END WL924
  PIN WL925
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 347.700 -1.950 347.900 ;
        RECT -3.750 347.100 -1.750 347.700 ;
        RECT -3.750 346.900 -1.950 347.100 ;
    END
  END WL925
  PIN WL926
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 345.450 -1.950 345.650 ;
        RECT -3.750 344.850 -1.750 345.450 ;
        RECT -3.750 344.650 -1.950 344.850 ;
    END
  END WL926
  PIN WL927
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 344.100 -1.950 344.300 ;
        RECT -3.750 343.500 -1.750 344.100 ;
        RECT -3.750 343.300 -1.950 343.500 ;
    END
  END WL927
  PIN WL928
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 341.850 -1.950 342.050 ;
        RECT -3.750 341.250 -1.750 341.850 ;
        RECT -3.750 341.050 -1.950 341.250 ;
    END
  END WL928
  PIN WL929
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 340.500 -1.950 340.700 ;
        RECT -3.750 339.900 -1.750 340.500 ;
        RECT -3.750 339.700 -1.950 339.900 ;
    END
  END WL929
  PIN WL930
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 338.250 -1.950 338.450 ;
        RECT -3.750 337.650 -1.750 338.250 ;
        RECT -3.750 337.450 -1.950 337.650 ;
    END
  END WL930
  PIN WL931
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 336.900 -1.950 337.100 ;
        RECT -3.750 336.300 -1.750 336.900 ;
        RECT -3.750 336.100 -1.950 336.300 ;
    END
  END WL931
  PIN WL932
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 334.650 -1.950 334.850 ;
        RECT -3.750 334.050 -1.750 334.650 ;
        RECT -3.750 333.850 -1.950 334.050 ;
    END
  END WL932
  PIN WL933
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 333.300 -1.950 333.500 ;
        RECT -3.750 332.700 -1.750 333.300 ;
        RECT -3.750 332.500 -1.950 332.700 ;
    END
  END WL933
  PIN WL934
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 331.050 -1.950 331.250 ;
        RECT -3.750 330.450 -1.750 331.050 ;
        RECT -3.750 330.250 -1.950 330.450 ;
    END
  END WL934
  PIN WL935
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 329.700 -1.950 329.900 ;
        RECT -3.750 329.100 -1.750 329.700 ;
        RECT -3.750 328.900 -1.950 329.100 ;
    END
  END WL935
  PIN WL936
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 327.450 -1.950 327.650 ;
        RECT -3.750 326.850 -1.750 327.450 ;
        RECT -3.750 326.650 -1.950 326.850 ;
    END
  END WL936
  PIN WL937
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 326.100 -1.950 326.300 ;
        RECT -3.750 325.500 -1.750 326.100 ;
        RECT -3.750 325.300 -1.950 325.500 ;
    END
  END WL937
  PIN WL938
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 323.850 -1.950 324.050 ;
        RECT -3.750 323.250 -1.750 323.850 ;
        RECT -3.750 323.050 -1.950 323.250 ;
    END
  END WL938
  PIN WL939
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 322.500 -1.950 322.700 ;
        RECT -3.750 321.900 -1.750 322.500 ;
        RECT -3.750 321.700 -1.950 321.900 ;
    END
  END WL939
  PIN WL940
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 320.250 -1.950 320.450 ;
        RECT -3.750 319.650 -1.750 320.250 ;
        RECT -3.750 319.450 -1.950 319.650 ;
    END
  END WL940
  PIN WL941
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 318.900 -1.950 319.100 ;
        RECT -3.750 318.300 -1.750 318.900 ;
        RECT -3.750 318.100 -1.950 318.300 ;
    END
  END WL941
  PIN WL942
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 316.650 -1.950 316.850 ;
        RECT -3.750 316.050 -1.750 316.650 ;
        RECT -3.750 315.850 -1.950 316.050 ;
    END
  END WL942
  PIN WL943
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 315.300 -1.950 315.500 ;
        RECT -3.750 314.700 -1.750 315.300 ;
        RECT -3.750 314.500 -1.950 314.700 ;
    END
  END WL943
  PIN WL944
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 313.050 -1.950 313.250 ;
        RECT -3.750 312.450 -1.750 313.050 ;
        RECT -3.750 312.250 -1.950 312.450 ;
    END
  END WL944
  PIN WL945
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 311.700 -1.950 311.900 ;
        RECT -3.750 311.100 -1.750 311.700 ;
        RECT -3.750 310.900 -1.950 311.100 ;
    END
  END WL945
  PIN WL946
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 309.450 -1.950 309.650 ;
        RECT -3.750 308.850 -1.750 309.450 ;
        RECT -3.750 308.650 -1.950 308.850 ;
    END
  END WL946
  PIN WL947
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 308.100 -1.950 308.300 ;
        RECT -3.750 307.500 -1.750 308.100 ;
        RECT -3.750 307.300 -1.950 307.500 ;
    END
  END WL947
  PIN WL948
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 305.850 -1.950 306.050 ;
        RECT -3.750 305.250 -1.750 305.850 ;
        RECT -3.750 305.050 -1.950 305.250 ;
    END
  END WL948
  PIN WL949
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 304.500 -1.950 304.700 ;
        RECT -3.750 303.900 -1.750 304.500 ;
        RECT -3.750 303.700 -1.950 303.900 ;
    END
  END WL949
  PIN WL950
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 302.250 -1.950 302.450 ;
        RECT -3.750 301.650 -1.750 302.250 ;
        RECT -3.750 301.450 -1.950 301.650 ;
    END
  END WL950
  PIN WL951
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 300.900 -1.950 301.100 ;
        RECT -3.750 300.300 -1.750 300.900 ;
        RECT -3.750 300.100 -1.950 300.300 ;
    END
  END WL951
  PIN WL952
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 298.650 -1.950 298.850 ;
        RECT -3.750 298.050 -1.750 298.650 ;
        RECT -3.750 297.850 -1.950 298.050 ;
    END
  END WL952
  PIN WL953
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 297.300 -1.950 297.500 ;
        RECT -3.750 296.700 -1.750 297.300 ;
        RECT -3.750 296.500 -1.950 296.700 ;
    END
  END WL953
  PIN WL954
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 295.050 -1.950 295.250 ;
        RECT -3.750 294.450 -1.750 295.050 ;
        RECT -3.750 294.250 -1.950 294.450 ;
    END
  END WL954
  PIN WL955
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 293.700 -1.950 293.900 ;
        RECT -3.750 293.100 -1.750 293.700 ;
        RECT -3.750 292.900 -1.950 293.100 ;
    END
  END WL955
  PIN WL956
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 291.450 -1.950 291.650 ;
        RECT -3.750 290.850 -1.750 291.450 ;
        RECT -3.750 290.650 -1.950 290.850 ;
    END
  END WL956
  PIN WL957
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 290.100 -1.950 290.300 ;
        RECT -3.750 289.500 -1.750 290.100 ;
        RECT -3.750 289.300 -1.950 289.500 ;
    END
  END WL957
  PIN WL958
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 287.850 -1.950 288.050 ;
        RECT -3.750 287.250 -1.750 287.850 ;
        RECT -3.750 287.050 -1.950 287.250 ;
    END
  END WL958
  PIN WL959
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 286.500 -1.950 286.700 ;
        RECT -3.750 285.900 -1.750 286.500 ;
        RECT -3.750 285.700 -1.950 285.900 ;
    END
  END WL959
  PIN WL960
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 284.250 -1.950 284.450 ;
        RECT -3.750 283.650 -1.750 284.250 ;
        RECT -3.750 283.450 -1.950 283.650 ;
    END
  END WL960
  PIN WL961
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 282.900 -1.950 283.100 ;
        RECT -3.750 282.300 -1.750 282.900 ;
        RECT -3.750 282.100 -1.950 282.300 ;
    END
  END WL961
  PIN WL962
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 280.650 -1.950 280.850 ;
        RECT -3.750 280.050 -1.750 280.650 ;
        RECT -3.750 279.850 -1.950 280.050 ;
    END
  END WL962
  PIN WL963
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 279.300 -1.950 279.500 ;
        RECT -3.750 278.700 -1.750 279.300 ;
        RECT -3.750 278.500 -1.950 278.700 ;
    END
  END WL963
  PIN WL964
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 277.050 -1.950 277.250 ;
        RECT -3.750 276.450 -1.750 277.050 ;
        RECT -3.750 276.250 -1.950 276.450 ;
    END
  END WL964
  PIN WL965
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 275.700 -1.950 275.900 ;
        RECT -3.750 275.100 -1.750 275.700 ;
        RECT -3.750 274.900 -1.950 275.100 ;
    END
  END WL965
  PIN WL966
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 273.450 -1.950 273.650 ;
        RECT -3.750 272.850 -1.750 273.450 ;
        RECT -3.750 272.650 -1.950 272.850 ;
    END
  END WL966
  PIN WL967
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 272.100 -1.950 272.300 ;
        RECT -3.750 271.500 -1.750 272.100 ;
        RECT -3.750 271.300 -1.950 271.500 ;
    END
  END WL967
  PIN WL968
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 269.850 -1.950 270.050 ;
        RECT -3.750 269.250 -1.750 269.850 ;
        RECT -3.750 269.050 -1.950 269.250 ;
    END
  END WL968
  PIN WL969
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 268.500 -1.950 268.700 ;
        RECT -3.750 267.900 -1.750 268.500 ;
        RECT -3.750 267.700 -1.950 267.900 ;
    END
  END WL969
  PIN WL970
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 266.250 -1.950 266.450 ;
        RECT -3.750 265.650 -1.750 266.250 ;
        RECT -3.750 265.450 -1.950 265.650 ;
    END
  END WL970
  PIN WL971
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 264.900 -1.950 265.100 ;
        RECT -3.750 264.300 -1.750 264.900 ;
        RECT -3.750 264.100 -1.950 264.300 ;
    END
  END WL971
  PIN WL972
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 262.650 -1.950 262.850 ;
        RECT -3.750 262.050 -1.750 262.650 ;
        RECT -3.750 261.850 -1.950 262.050 ;
    END
  END WL972
  PIN WL973
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 261.300 -1.950 261.500 ;
        RECT -3.750 260.700 -1.750 261.300 ;
        RECT -3.750 260.500 -1.950 260.700 ;
    END
  END WL973
  PIN WL974
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 259.050 -1.950 259.250 ;
        RECT -3.750 258.450 -1.750 259.050 ;
        RECT -3.750 258.250 -1.950 258.450 ;
    END
  END WL974
  PIN WL975
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 257.700 -1.950 257.900 ;
        RECT -3.750 257.100 -1.750 257.700 ;
        RECT -3.750 256.900 -1.950 257.100 ;
    END
  END WL975
  PIN WL976
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 255.450 -1.950 255.650 ;
        RECT -3.750 254.850 -1.750 255.450 ;
        RECT -3.750 254.650 -1.950 254.850 ;
    END
  END WL976
  PIN WL977
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 254.100 -1.950 254.300 ;
        RECT -3.750 253.500 -1.750 254.100 ;
        RECT -3.750 253.300 -1.950 253.500 ;
    END
  END WL977
  PIN WL978
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 251.850 -1.950 252.050 ;
        RECT -3.750 251.250 -1.750 251.850 ;
        RECT -3.750 251.050 -1.950 251.250 ;
    END
  END WL978
  PIN WL979
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 250.500 -1.950 250.700 ;
        RECT -3.750 249.900 -1.750 250.500 ;
        RECT -3.750 249.700 -1.950 249.900 ;
    END
  END WL979
  PIN WL980
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 248.250 -1.950 248.450 ;
        RECT -3.750 247.650 -1.750 248.250 ;
        RECT -3.750 247.450 -1.950 247.650 ;
    END
  END WL980
  PIN WL981
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 246.900 -1.950 247.100 ;
        RECT -3.750 246.300 -1.750 246.900 ;
        RECT -3.750 246.100 -1.950 246.300 ;
    END
  END WL981
  PIN WL982
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 244.650 -1.950 244.850 ;
        RECT -3.750 244.050 -1.750 244.650 ;
        RECT -3.750 243.850 -1.950 244.050 ;
    END
  END WL982
  PIN WL983
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 243.300 -1.950 243.500 ;
        RECT -3.750 242.700 -1.750 243.300 ;
        RECT -3.750 242.500 -1.950 242.700 ;
    END
  END WL983
  PIN WL984
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 241.050 -1.950 241.250 ;
        RECT -3.750 240.450 -1.750 241.050 ;
        RECT -3.750 240.250 -1.950 240.450 ;
    END
  END WL984
  PIN WL985
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 239.700 -1.950 239.900 ;
        RECT -3.750 239.100 -1.750 239.700 ;
        RECT -3.750 238.900 -1.950 239.100 ;
    END
  END WL985
  PIN WL986
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 237.450 -1.950 237.650 ;
        RECT -3.750 236.850 -1.750 237.450 ;
        RECT -3.750 236.650 -1.950 236.850 ;
    END
  END WL986
  PIN WL987
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 236.100 -1.950 236.300 ;
        RECT -3.750 235.500 -1.750 236.100 ;
        RECT -3.750 235.300 -1.950 235.500 ;
    END
  END WL987
  PIN WL988
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 233.850 -1.950 234.050 ;
        RECT -3.750 233.250 -1.750 233.850 ;
        RECT -3.750 233.050 -1.950 233.250 ;
    END
  END WL988
  PIN WL989
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 232.500 -1.950 232.700 ;
        RECT -3.750 231.900 -1.750 232.500 ;
        RECT -3.750 231.700 -1.950 231.900 ;
    END
  END WL989
  PIN WL990
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 230.250 -1.950 230.450 ;
        RECT -3.750 229.650 -1.750 230.250 ;
        RECT -3.750 229.450 -1.950 229.650 ;
    END
  END WL990
  PIN WL991
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 228.900 -1.950 229.100 ;
        RECT -3.750 228.300 -1.750 228.900 ;
        RECT -3.750 228.100 -1.950 228.300 ;
    END
  END WL991
  PIN WL992
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 226.650 -1.950 226.850 ;
        RECT -3.750 226.050 -1.750 226.650 ;
        RECT -3.750 225.850 -1.950 226.050 ;
    END
  END WL992
  PIN WL993
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 225.300 -1.950 225.500 ;
        RECT -3.750 224.700 -1.750 225.300 ;
        RECT -3.750 224.500 -1.950 224.700 ;
    END
  END WL993
  PIN WL994
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 222.500 -1.950 222.700 ;
        RECT -3.750 221.900 -1.750 222.500 ;
        RECT -3.750 221.700 -1.950 221.900 ;
    END
  END WL994
  PIN WL995
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 221.150 -1.950 221.350 ;
        RECT -3.750 220.550 -1.750 221.150 ;
        RECT -3.750 220.350 -1.950 220.550 ;
    END
  END WL995
  PIN WL996
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 218.900 -1.950 219.100 ;
        RECT -3.750 218.300 -1.750 218.900 ;
        RECT -3.750 218.100 -1.950 218.300 ;
    END
  END WL996
  PIN WL997
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 217.550 -1.950 217.750 ;
        RECT -3.750 216.950 -1.750 217.550 ;
        RECT -3.750 216.750 -1.950 216.950 ;
    END
  END WL997
  PIN WL998
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 215.300 -1.950 215.500 ;
        RECT -3.750 214.700 -1.750 215.300 ;
        RECT -3.750 214.500 -1.950 214.700 ;
    END
  END WL998
  PIN WL999
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 213.950 -1.950 214.150 ;
        RECT -3.750 213.350 -1.750 213.950 ;
        RECT -3.750 213.150 -1.950 213.350 ;
    END
  END WL999
  PIN WL1000
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 211.700 -1.950 211.900 ;
        RECT -3.750 211.100 -1.750 211.700 ;
        RECT -3.750 210.900 -1.950 211.100 ;
    END
  END WL1000
  PIN WL1001
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 210.350 -1.950 210.550 ;
        RECT -3.750 209.750 -1.750 210.350 ;
        RECT -3.750 209.550 -1.950 209.750 ;
    END
  END WL1001
  PIN WL1002
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 208.100 -1.950 208.300 ;
        RECT -3.750 207.500 -1.750 208.100 ;
        RECT -3.750 207.300 -1.950 207.500 ;
    END
  END WL1002
  PIN WL1003
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 206.750 -1.950 206.950 ;
        RECT -3.750 206.150 -1.750 206.750 ;
        RECT -3.750 205.950 -1.950 206.150 ;
    END
  END WL1003
  PIN WL1004
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 204.500 -1.950 204.700 ;
        RECT -3.750 203.900 -1.750 204.500 ;
        RECT -3.750 203.700 -1.950 203.900 ;
    END
  END WL1004
  PIN WL1005
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 203.150 -1.950 203.350 ;
        RECT -3.750 202.550 -1.750 203.150 ;
        RECT -3.750 202.350 -1.950 202.550 ;
    END
  END WL1005
  PIN WL1006
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 200.900 -1.950 201.100 ;
        RECT -3.750 200.300 -1.750 200.900 ;
        RECT -3.750 200.100 -1.950 200.300 ;
    END
  END WL1006
  PIN WL1007
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 199.550 -1.950 199.750 ;
        RECT -3.750 198.950 -1.750 199.550 ;
        RECT -3.750 198.750 -1.950 198.950 ;
    END
  END WL1007
  PIN WL1008
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 197.300 -1.950 197.500 ;
        RECT -3.750 196.700 -1.750 197.300 ;
        RECT -3.750 196.500 -1.950 196.700 ;
    END
  END WL1008
  PIN WL1009
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 195.950 -1.950 196.150 ;
        RECT -3.750 195.350 -1.750 195.950 ;
        RECT -3.750 195.150 -1.950 195.350 ;
    END
  END WL1009
  PIN WL1010
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 193.700 -1.950 193.900 ;
        RECT -3.750 193.100 -1.750 193.700 ;
        RECT -3.750 192.900 -1.950 193.100 ;
    END
  END WL1010
  PIN WL1011
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 192.350 -1.950 192.550 ;
        RECT -3.750 191.750 -1.750 192.350 ;
        RECT -3.750 191.550 -1.950 191.750 ;
    END
  END WL1011
  PIN WL1012
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 190.100 -1.950 190.300 ;
        RECT -3.750 189.500 -1.750 190.100 ;
        RECT -3.750 189.300 -1.950 189.500 ;
    END
  END WL1012
  PIN WL1013
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 188.750 -1.950 188.950 ;
        RECT -3.750 188.150 -1.750 188.750 ;
        RECT -3.750 187.950 -1.950 188.150 ;
    END
  END WL1013
  PIN WL1014
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 186.500 -1.950 186.700 ;
        RECT -3.750 185.900 -1.750 186.500 ;
        RECT -3.750 185.700 -1.950 185.900 ;
    END
  END WL1014
  PIN WL1015
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 185.150 -1.950 185.350 ;
        RECT -3.750 184.550 -1.750 185.150 ;
        RECT -3.750 184.350 -1.950 184.550 ;
    END
  END WL1015
  PIN WL1016
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 182.900 -1.950 183.100 ;
        RECT -3.750 182.300 -1.750 182.900 ;
        RECT -3.750 182.100 -1.950 182.300 ;
    END
  END WL1016
  PIN WL1017
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 181.550 -1.950 181.750 ;
        RECT -3.750 180.950 -1.750 181.550 ;
        RECT -3.750 180.750 -1.950 180.950 ;
    END
  END WL1017
  PIN WL1018
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 179.300 -1.950 179.500 ;
        RECT -3.750 178.700 -1.750 179.300 ;
        RECT -3.750 178.500 -1.950 178.700 ;
    END
  END WL1018
  PIN WL1019
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 177.950 -1.950 178.150 ;
        RECT -3.750 177.350 -1.750 177.950 ;
        RECT -3.750 177.150 -1.950 177.350 ;
    END
  END WL1019
  PIN WL1020
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 175.700 -1.950 175.900 ;
        RECT -3.750 175.100 -1.750 175.700 ;
        RECT -3.750 174.900 -1.950 175.100 ;
    END
  END WL1020
  PIN WL1021
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 174.350 -1.950 174.550 ;
        RECT -3.750 173.750 -1.750 174.350 ;
        RECT -3.750 173.550 -1.950 173.750 ;
    END
  END WL1021
  PIN WL1022
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 172.100 -1.950 172.300 ;
        RECT -3.750 171.500 -1.750 172.100 ;
        RECT -3.750 171.300 -1.950 171.500 ;
    END
  END WL1022
  PIN WL1023
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -3.750 170.750 -1.950 170.950 ;
        RECT -3.750 170.150 -1.750 170.750 ;
        RECT -3.750 169.950 -1.950 170.150 ;
    END
  END WL1023
  OBS
      LAYER li1 ;
        RECT 13.000 29.150 246.980 2022.680 ;
      LAYER met1 ;
        RECT 7.250 19.900 247.640 2023.350 ;
      LAYER met2 ;
        RECT -1.750 19.900 257.250 2031.600 ;
      LAYER met3 ;
        RECT -1.950 36.000 257.250 2028.600 ;
      LAYER met4 ;
        RECT 92.500 86.500 220.900 89.100 ;
  END
END truncation_SRAM
END LIBRARY

