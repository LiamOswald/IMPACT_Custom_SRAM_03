magic
tech sky130B
magscale 1 2
timestamp 1713986195
<< metal1 >>
rect 494790 700272 494796 700324
rect 494848 700312 494854 700324
rect 512086 700312 512092 700324
rect 494848 700284 512092 700312
rect 494848 700272 494854 700284
rect 512086 700272 512092 700284
rect 512144 700272 512150 700324
rect 502242 1300 502248 1352
rect 502300 1340 502306 1352
rect 511994 1340 512000 1352
rect 502300 1312 512000 1340
rect 502300 1300 502306 1312
rect 511994 1300 512000 1312
rect 512052 1300 512058 1352
rect 3602 1232 3608 1284
rect 3660 1272 3666 1284
rect 155954 1272 155960 1284
rect 3660 1244 155960 1272
rect 3660 1232 3666 1244
rect 155954 1232 155960 1244
rect 156012 1232 156018 1284
rect 368382 1232 368388 1284
rect 368440 1272 368446 1284
rect 559650 1272 559656 1284
rect 368440 1244 559656 1272
rect 368440 1232 368446 1244
rect 559650 1232 559656 1244
rect 559708 1232 559714 1284
rect 3510 1164 3516 1216
rect 3568 1204 3574 1216
rect 136634 1204 136640 1216
rect 3568 1176 136640 1204
rect 3568 1164 3574 1176
rect 136634 1164 136640 1176
rect 136692 1164 136698 1216
rect 406470 1164 406476 1216
rect 406528 1204 406534 1216
rect 580350 1204 580356 1216
rect 406528 1176 580356 1204
rect 406528 1164 406534 1176
rect 580350 1164 580356 1176
rect 580408 1164 580414 1216
rect 3418 1096 3424 1148
rect 3476 1136 3482 1148
rect 117406 1136 117412 1148
rect 3476 1108 117412 1136
rect 3476 1096 3482 1108
rect 117406 1096 117412 1108
rect 117464 1096 117470 1148
rect 445662 1096 445668 1148
rect 445720 1136 445726 1148
rect 580442 1136 580448 1148
rect 445720 1108 580448 1136
rect 445720 1096 445726 1108
rect 580442 1096 580448 1108
rect 580500 1096 580506 1148
rect 387702 1028 387708 1080
rect 387760 1068 387766 1080
rect 512086 1068 512092 1080
rect 387760 1040 512092 1068
rect 387760 1028 387766 1040
rect 512086 1028 512092 1040
rect 512144 1028 512150 1080
rect 483382 960 483388 1012
rect 483440 1000 483446 1012
rect 511350 1000 511356 1012
rect 483440 972 511356 1000
rect 483440 960 483446 972
rect 511350 960 511356 972
rect 511408 960 511414 1012
rect 21910 892 21916 944
rect 21968 932 21974 944
rect 580258 932 580264 944
rect 21968 904 580264 932
rect 21968 892 21974 904
rect 580258 892 580264 904
rect 580316 892 580322 944
<< via1 >>
rect 494796 700272 494848 700324
rect 512092 700272 512144 700324
rect 502248 1300 502300 1352
rect 512000 1300 512052 1352
rect 3608 1232 3660 1284
rect 155960 1232 156012 1284
rect 368388 1232 368440 1284
rect 559656 1232 559708 1284
rect 3516 1164 3568 1216
rect 136640 1164 136692 1216
rect 406476 1164 406528 1216
rect 580356 1164 580408 1216
rect 3424 1096 3476 1148
rect 117412 1096 117464 1148
rect 445668 1096 445720 1148
rect 580448 1096 580500 1148
rect 387708 1028 387760 1080
rect 512092 1028 512144 1080
rect 483388 960 483440 1012
rect 511356 960 511408 1012
rect 21916 892 21968 944
rect 580264 892 580316 944
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 9586 700904 9642 700913
rect 9586 700839 9642 700848
rect 9494 700768 9550 700777
rect 9494 700703 9550 700712
rect 9310 700632 9366 700641
rect 9310 700567 9366 700576
rect 9324 502761 9352 700567
rect 9402 700496 9458 700505
rect 9402 700431 9458 700440
rect 9310 502752 9366 502761
rect 9310 502687 9366 502696
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2962 71632 3018 71641
rect 2962 71567 3018 71576
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 2792 921 2820 32399
rect 2976 1057 3004 71567
rect 3160 1329 3188 110599
rect 3146 1320 3202 1329
rect 3146 1255 3202 1264
rect 3344 1193 3372 162823
rect 3330 1184 3386 1193
rect 3436 1154 3464 475623
rect 9416 436121 9444 700431
rect 9402 436112 9458 436121
rect 9402 436047 9458 436056
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 1222 3556 423535
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3620 1290 3648 371311
rect 9508 369481 9536 700703
rect 9494 369472 9550 369481
rect 9494 369407 9550 369416
rect 3698 319288 3754 319297
rect 3698 319223 3754 319232
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 3330 1119 3386 1128
rect 3424 1148 3476 1154
rect 3424 1090 3476 1096
rect 2962 1048 3018 1057
rect 2962 983 3018 992
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 3712 513 3740 319223
rect 9600 302841 9628 700839
rect 56796 700369 56824 703520
rect 121656 700641 121684 703520
rect 186516 700641 186544 703520
rect 235184 700913 235212 703520
rect 235170 700904 235226 700913
rect 235170 700839 235226 700848
rect 262034 700904 262090 700913
rect 262034 700839 262090 700848
rect 121642 700632 121698 700641
rect 121642 700567 121698 700576
rect 186502 700632 186558 700641
rect 186502 700567 186558 700576
rect 56782 700360 56838 700369
rect 56782 700295 56838 700304
rect 262048 603242 262076 700839
rect 300136 700777 300164 703520
rect 300122 700768 300178 700777
rect 300122 700703 300178 700712
rect 364996 700505 365024 703520
rect 429856 700913 429884 703520
rect 429842 700904 429898 700913
rect 429842 700839 429898 700848
rect 364982 700496 365038 700505
rect 364982 700431 365038 700440
rect 494808 700330 494836 703520
rect 511998 700632 512054 700641
rect 511998 700567 512054 700576
rect 511354 700360 511410 700369
rect 494796 700324 494848 700330
rect 511354 700295 511410 700304
rect 494796 700266 494848 700272
rect 262002 603214 262076 603242
rect 262002 602956 262030 603214
rect 9586 302832 9642 302841
rect 9586 302767 9642 302776
rect 3882 267200 3938 267209
rect 3882 267135 3938 267144
rect 3896 649 3924 267135
rect 4066 214976 4122 214985
rect 4066 214911 4122 214920
rect 4080 785 4108 214911
rect 425380 3088 425436 3097
rect 21620 3046 21956 3074
rect 21928 950 21956 3046
rect 40512 3046 40848 3074
rect 59740 3046 60076 3074
rect 79304 3046 79548 3074
rect 98532 3046 98868 3074
rect 21916 944 21968 950
rect 40512 921 40540 3046
rect 59740 1057 59768 3046
rect 59726 1048 59782 1057
rect 59726 983 59782 992
rect 21916 886 21968 892
rect 40498 912 40554 921
rect 40498 847 40554 856
rect 4066 776 4122 785
rect 4066 711 4122 720
rect 3882 640 3938 649
rect 3882 575 3938 584
rect 3698 504 3754 513
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3698 439 3754 448
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79520 377 79548 3046
rect 98840 921 98868 3046
rect 117424 3046 117760 3074
rect 136652 3046 136988 3074
rect 155972 3046 156216 3074
rect 175292 3046 175444 3074
rect 194612 3046 194672 3074
rect 213564 3046 213900 3074
rect 232792 3046 233128 3074
rect 252020 3046 252356 3074
rect 271584 3046 271828 3074
rect 290812 3046 291148 3074
rect 310040 3046 310376 3074
rect 329268 3046 329604 3074
rect 348496 3046 348832 3074
rect 367724 3046 368060 3074
rect 117424 1154 117452 3046
rect 136652 1222 136680 3046
rect 155972 1290 156000 3046
rect 155960 1284 156012 1290
rect 155960 1226 156012 1232
rect 136640 1216 136692 1222
rect 136640 1158 136692 1164
rect 117412 1148 117464 1154
rect 117412 1090 117464 1096
rect 98826 912 98882 921
rect 98826 847 98882 856
rect 175292 513 175320 3046
rect 194612 649 194640 3046
rect 213564 785 213592 3046
rect 232792 1193 232820 3046
rect 252020 1329 252048 3046
rect 271800 1329 271828 3046
rect 252006 1320 252062 1329
rect 252006 1255 252062 1264
rect 271786 1320 271842 1329
rect 271786 1255 271842 1264
rect 291120 1193 291148 3046
rect 232778 1184 232834 1193
rect 232778 1119 232834 1128
rect 291106 1184 291162 1193
rect 291106 1119 291162 1128
rect 310348 785 310376 3046
rect 213550 776 213606 785
rect 213550 711 213606 720
rect 310334 776 310390 785
rect 310334 711 310390 720
rect 329576 649 329604 3046
rect 348804 1057 348832 3046
rect 348790 1048 348846 1057
rect 348790 983 348846 992
rect 194598 640 194654 649
rect 194598 575 194654 584
rect 329562 640 329618 649
rect 329562 575 329618 584
rect 368032 513 368060 3046
rect 386892 3046 386952 3074
rect 406180 3046 406516 3074
rect 368388 1284 368440 1290
rect 368388 1226 368440 1232
rect 175278 504 175334 513
rect 79506 368 79562 377
rect 79506 303 79562 312
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 368018 504 368074 513
rect 175278 439 175334 448
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368018 439 368074 448
rect 368174 -960 368286 480
rect 368400 377 368428 1226
rect 368386 368 368442 377
rect 368386 303 368442 312
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386892 377 386920 3046
rect 406488 1222 406516 3046
rect 444636 3046 444880 3074
rect 425380 3023 425436 3032
rect 406476 1216 406528 1222
rect 406476 1158 406528 1164
rect 387708 1080 387760 1086
rect 387708 1022 387760 1028
rect 387720 921 387748 1022
rect 387706 912 387762 921
rect 387706 847 387762 856
rect 386878 368 386934 377
rect 386878 303 386934 312
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444852 105 444880 3046
rect 463850 2961 463878 3060
rect 483092 3046 483428 3074
rect 463836 2952 463892 2961
rect 463836 2887 463892 2896
rect 445668 1148 445720 1154
rect 445668 1090 445720 1096
rect 444838 96 444894 105
rect 444838 31 444894 40
rect 444994 -960 445106 480
rect 445680 377 445708 1090
rect 483400 1018 483428 3046
rect 502260 3046 502320 3074
rect 502260 1358 502288 3046
rect 502248 1352 502300 1358
rect 502248 1294 502300 1300
rect 511368 1018 511396 700295
rect 512012 1358 512040 700567
rect 512092 700324 512144 700330
rect 512092 700266 512144 700272
rect 512000 1352 512052 1358
rect 512000 1294 512052 1300
rect 512104 1086 512132 700266
rect 514022 347712 514078 347721
rect 514022 347647 514078 347656
rect 514036 232393 514064 347647
rect 514206 287872 514262 287881
rect 514206 287807 514262 287816
rect 514022 232384 514078 232393
rect 514022 232319 514078 232328
rect 514114 228032 514170 228041
rect 514114 227967 514170 227976
rect 514022 198112 514078 198121
rect 514022 198047 514078 198056
rect 514036 33153 514064 198047
rect 514128 73001 514156 227967
rect 514220 152697 514248 287807
rect 514206 152688 514262 152697
rect 514206 152623 514262 152632
rect 514114 72992 514170 73001
rect 514114 72927 514170 72936
rect 514022 33144 514078 33153
rect 514022 33079 514078 33088
rect 559668 1290 559696 703520
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 579816 1329 579844 258839
rect 579802 1320 579858 1329
rect 559656 1284 559708 1290
rect 579802 1255 579858 1264
rect 559656 1226 559708 1232
rect 580000 1193 580028 312015
rect 579986 1184 580042 1193
rect 579986 1119 580042 1128
rect 512092 1080 512144 1086
rect 512092 1022 512144 1028
rect 483388 1012 483440 1018
rect 483388 954 483440 960
rect 511356 1012 511408 1018
rect 511356 954 511408 960
rect 580184 785 580212 365055
rect 580276 950 580304 670647
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580368 1222 580396 630799
rect 580446 577688 580502 577697
rect 580446 577623 580502 577632
rect 580356 1216 580408 1222
rect 580356 1158 580408 1164
rect 580460 1154 580488 577623
rect 580538 524512 580594 524521
rect 580538 524447 580594 524456
rect 580448 1148 580500 1154
rect 580448 1090 580500 1096
rect 580264 944 580316 950
rect 580264 886 580316 892
rect 580170 776 580226 785
rect 580170 711 580226 720
rect 580552 513 580580 524447
rect 580722 471472 580778 471481
rect 580722 471407 580778 471416
rect 580736 1057 580764 471407
rect 580906 418296 580962 418305
rect 580906 418231 580962 418240
rect 580722 1048 580778 1057
rect 580722 983 580778 992
rect 580920 649 580948 418231
rect 580998 3088 581054 3097
rect 580998 3023 581054 3032
rect 580906 640 580962 649
rect 580906 575 580962 584
rect 580538 504 580594 513
rect 445666 368 445722 377
rect 445666 303 445722 312
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 581012 480 581040 3023
rect 583390 2952 583446 2961
rect 583390 2887 583446 2896
rect 583404 480 583432 2887
rect 580538 439 580594 448
rect 580970 -960 581082 480
rect 581826 96 581882 105
rect 582166 82 582278 480
rect 581882 54 582278 82
rect 581826 31 581882 40
rect 582166 -960 582278 54
rect 583362 -960 583474 480
<< via2 >>
rect 9586 700848 9642 700904
rect 9494 700712 9550 700768
rect 9310 700576 9366 700632
rect 9402 700440 9458 700496
rect 9310 502696 9366 502752
rect 3422 475632 3478 475688
rect 3330 162832 3386 162888
rect 3146 110608 3202 110664
rect 2962 71576 3018 71632
rect 2778 32408 2834 32464
rect 3146 1264 3202 1320
rect 3330 1128 3386 1184
rect 9402 436056 9458 436112
rect 3514 423544 3570 423600
rect 3606 371320 3662 371376
rect 9494 369416 9550 369472
rect 3698 319232 3754 319288
rect 2962 992 3018 1048
rect 2778 856 2834 912
rect 235170 700848 235226 700904
rect 262034 700848 262090 700904
rect 121642 700576 121698 700632
rect 186502 700576 186558 700632
rect 56782 700304 56838 700360
rect 300122 700712 300178 700768
rect 429842 700848 429898 700904
rect 364982 700440 365038 700496
rect 511998 700576 512054 700632
rect 511354 700304 511410 700360
rect 9586 302776 9642 302832
rect 3882 267144 3938 267200
rect 4066 214920 4122 214976
rect 59726 992 59782 1048
rect 40498 856 40554 912
rect 4066 720 4122 776
rect 3882 584 3938 640
rect 3698 448 3754 504
rect 98826 856 98882 912
rect 252006 1264 252062 1320
rect 271786 1264 271842 1320
rect 232778 1128 232834 1184
rect 291106 1128 291162 1184
rect 213550 720 213606 776
rect 310334 720 310390 776
rect 348790 992 348846 1048
rect 194598 584 194654 640
rect 329562 584 329618 640
rect 79506 312 79562 368
rect 175278 448 175334 504
rect 368018 448 368074 504
rect 368386 312 368442 368
rect 425380 3032 425436 3088
rect 387706 856 387762 912
rect 386878 312 386934 368
rect 463836 2896 463892 2952
rect 444838 40 444894 96
rect 514022 347656 514078 347712
rect 514206 287816 514262 287872
rect 514022 232328 514078 232384
rect 514114 227976 514170 228032
rect 514022 198056 514078 198112
rect 514206 152632 514262 152688
rect 514114 72936 514170 72992
rect 514022 33088 514078 33144
rect 580262 670656 580318 670712
rect 580170 365064 580226 365120
rect 579986 312024 580042 312080
rect 579802 258848 579858 258904
rect 579802 1264 579858 1320
rect 579986 1128 580042 1184
rect 580354 630808 580410 630864
rect 580446 577632 580502 577688
rect 580538 524456 580594 524512
rect 580170 720 580226 776
rect 580722 471416 580778 471472
rect 580906 418240 580962 418296
rect 580722 992 580778 1048
rect 580998 3032 581054 3088
rect 580906 584 580962 640
rect 445666 312 445722 368
rect 580538 448 580594 504
rect 583390 2896 583446 2952
rect 581826 40 581882 96
<< metal3 >>
rect 9581 700906 9647 700909
rect 235165 700906 235231 700909
rect 9581 700904 235231 700906
rect 9581 700848 9586 700904
rect 9642 700848 235170 700904
rect 235226 700848 235231 700904
rect 9581 700846 235231 700848
rect 9581 700843 9647 700846
rect 235165 700843 235231 700846
rect 262029 700906 262095 700909
rect 429837 700906 429903 700909
rect 262029 700904 429903 700906
rect 262029 700848 262034 700904
rect 262090 700848 429842 700904
rect 429898 700848 429903 700904
rect 262029 700846 429903 700848
rect 262029 700843 262095 700846
rect 429837 700843 429903 700846
rect 9489 700770 9555 700773
rect 300117 700770 300183 700773
rect 9489 700768 300183 700770
rect 9489 700712 9494 700768
rect 9550 700712 300122 700768
rect 300178 700712 300183 700768
rect 9489 700710 300183 700712
rect 9489 700707 9555 700710
rect 300117 700707 300183 700710
rect 9305 700634 9371 700637
rect 121637 700634 121703 700637
rect 9305 700632 121703 700634
rect 9305 700576 9310 700632
rect 9366 700576 121642 700632
rect 121698 700576 121703 700632
rect 9305 700574 121703 700576
rect 9305 700571 9371 700574
rect 121637 700571 121703 700574
rect 186497 700634 186563 700637
rect 511993 700634 512059 700637
rect 186497 700632 512059 700634
rect 186497 700576 186502 700632
rect 186558 700576 511998 700632
rect 512054 700576 512059 700632
rect 186497 700574 512059 700576
rect 186497 700571 186563 700574
rect 511993 700571 512059 700574
rect 9397 700498 9463 700501
rect 364977 700498 365043 700501
rect 9397 700496 365043 700498
rect 9397 700440 9402 700496
rect 9458 700440 364982 700496
rect 365038 700440 365043 700496
rect 9397 700438 365043 700440
rect 9397 700435 9463 700438
rect 364977 700435 365043 700438
rect 56777 700362 56843 700365
rect 511349 700362 511415 700365
rect 56777 700360 511415 700362
rect 56777 700304 56782 700360
rect 56838 700304 511354 700360
rect 511410 700304 511415 700360
rect 56777 700302 511415 700304
rect 56777 700299 56843 700302
rect 511349 700299 511415 700302
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3550 684314 3556 684316
rect -960 684254 3556 684314
rect -960 684164 480 684254
rect 3550 684252 3556 684254
rect 3620 684252 3626 684316
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 514150 643996 514156 644060
rect 514220 644058 514226 644060
rect 583520 644058 584960 644148
rect 514220 643998 584960 644058
rect 514220 643996 514226 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3918 632090 3924 632092
rect -960 632030 3924 632090
rect -960 631940 480 632030
rect 3918 632028 3924 632030
rect 3988 632028 3994 632092
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 583520 630716 584960 630806
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect 12014 602244 12020 602308
rect 12084 602306 12090 602308
rect 580206 602306 580212 602308
rect 12084 602246 580212 602306
rect 12084 602244 12090 602246
rect 580206 602244 580212 602246
rect 580276 602244 580282 602308
rect -960 592908 480 593148
rect 580390 590956 580396 591020
rect 580460 591018 580466 591020
rect 583520 591018 584960 591108
rect 580460 590958 584960 591018
rect 580460 590956 580466 590958
rect 583520 590868 584960 590958
rect 514150 587074 514156 587076
rect 511796 587014 514156 587074
rect 514150 587012 514156 587014
rect 514220 587012 514226 587076
rect -960 580002 480 580092
rect 3366 580002 3372 580004
rect -960 579942 3372 580002
rect -960 579852 480 579942
rect 3366 579940 3372 579942
rect 3436 579940 3442 580004
rect 580441 577690 580507 577693
rect 583520 577690 584960 577780
rect 580441 577688 584960 577690
rect 580441 577632 580446 577688
rect 580502 577632 584960 577688
rect 580441 577630 584960 577632
rect 580441 577627 580507 577630
rect 583520 577540 584960 577630
rect 12014 569332 12020 569396
rect 12084 569332 12090 569396
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect 580390 557154 580396 557156
rect 511796 557094 580396 557154
rect 580390 557092 580396 557094
rect 580460 557092 580466 557156
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 514150 537780 514156 537844
rect 514220 537842 514226 537844
rect 583520 537842 584960 537932
rect 514220 537782 584960 537842
rect 514220 537780 514226 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3734 527914 3740 527916
rect -960 527854 3740 527914
rect -960 527764 480 527854
rect 3734 527852 3740 527854
rect 3804 527852 3810 527916
rect 514150 527234 514156 527236
rect 511796 527174 514156 527234
rect 514150 527172 514156 527174
rect 514220 527172 514226 527236
rect 580533 524514 580599 524517
rect 583520 524514 584960 524604
rect 580533 524512 584960 524514
rect 580533 524456 580538 524512
rect 580594 524456 584960 524512
rect 580533 524454 584960 524456
rect 580533 524451 580599 524454
rect 583520 524364 584960 524454
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect 9305 502754 9371 502757
rect 9305 502752 12052 502754
rect 9305 502696 9310 502752
rect 9366 502696 12052 502752
rect 9305 502694 12052 502696
rect 9305 502691 9371 502694
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 514150 497314 514156 497316
rect 511796 497254 514156 497314
rect 514150 497252 514156 497254
rect 514220 497252 514226 497316
rect -960 488596 480 488836
rect 514150 484604 514156 484668
rect 514220 484666 514226 484668
rect 583520 484666 584960 484756
rect 514220 484606 584960 484666
rect 514220 484604 514226 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580717 471474 580783 471477
rect 583520 471474 584960 471564
rect 580717 471472 584960 471474
rect 580717 471416 580722 471472
rect 580778 471416 584960 471472
rect 580717 471414 584960 471416
rect 580717 471411 580783 471414
rect 583520 471324 584960 471414
rect 514334 467394 514340 467396
rect 511796 467334 514340 467394
rect 514334 467332 514340 467334
rect 514404 467332 514410 467396
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect 514150 437474 514156 437476
rect 511796 437414 514156 437474
rect 514150 437412 514156 437414
rect 514220 437412 514226 437476
rect -960 436508 480 436748
rect 9397 436114 9463 436117
rect 9397 436112 12052 436114
rect 9397 436056 9402 436112
rect 9458 436056 12052 436112
rect 9397 436054 12052 436056
rect 9397 436051 9463 436054
rect 514334 431564 514340 431628
rect 514404 431626 514410 431628
rect 583520 431626 584960 431716
rect 514404 431566 584960 431626
rect 514404 431564 514410 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580901 418298 580967 418301
rect 583520 418298 584960 418388
rect 580901 418296 584960 418298
rect 580901 418240 580906 418296
rect 580962 418240 584960 418296
rect 580901 418238 584960 418240
rect 580901 418235 580967 418238
rect 583520 418148 584960 418238
rect -960 410396 480 410636
rect 514334 407554 514340 407556
rect 511796 407494 514340 407554
rect 514334 407492 514340 407494
rect 514404 407492 514410 407556
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 514150 378388 514156 378452
rect 514220 378450 514226 378452
rect 583520 378450 584960 378540
rect 514220 378390 584960 378450
rect 514220 378388 514226 378390
rect 583520 378300 584960 378390
rect 514150 377634 514156 377636
rect 511796 377574 514156 377634
rect 514150 377572 514156 377574
rect 514220 377572 514226 377636
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 9489 369474 9555 369477
rect 9489 369472 12052 369474
rect 9489 369416 9494 369472
rect 9550 369416 12052 369472
rect 9489 369414 12052 369416
rect 9489 369411 9555 369414
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect 514017 347714 514083 347717
rect 511796 347712 514083 347714
rect 511796 347656 514022 347712
rect 514078 347656 514083 347712
rect 511796 347654 514083 347656
rect 514017 347651 514083 347654
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 514334 325212 514340 325276
rect 514404 325274 514410 325276
rect 583520 325274 584960 325364
rect 514404 325214 584960 325274
rect 514404 325212 514410 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3693 319290 3759 319293
rect -960 319288 3759 319290
rect -960 319232 3698 319288
rect 3754 319232 3759 319288
rect -960 319230 3759 319232
rect -960 319140 480 319230
rect 3693 319227 3759 319230
rect 514334 317794 514340 317796
rect 511796 317734 514340 317794
rect 514334 317732 514340 317734
rect 514404 317732 514410 317796
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306084 480 306324
rect 9581 302834 9647 302837
rect 9581 302832 12052 302834
rect 9581 302776 9586 302832
rect 9642 302776 12052 302832
rect 9581 302774 12052 302776
rect 9581 302771 9647 302774
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 514201 287874 514267 287877
rect 511796 287872 514267 287874
rect 511796 287816 514206 287872
rect 514262 287816 514267 287872
rect 511796 287814 514267 287816
rect 514201 287811 514267 287814
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 514150 272172 514156 272236
rect 514220 272234 514226 272236
rect 583520 272234 584960 272324
rect 514220 272174 584960 272234
rect 514220 272172 514226 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3877 267202 3943 267205
rect -960 267200 3943 267202
rect -960 267144 3882 267200
rect 3938 267144 3943 267200
rect -960 267142 3943 267144
rect -960 267052 480 267142
rect 3877 267139 3943 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect 514150 257954 514156 257956
rect 511796 257894 514156 257954
rect 514150 257892 514156 257894
rect 514220 257892 514226 257956
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 3918 236132 3924 236196
rect 3988 236194 3994 236196
rect 3988 236134 12052 236194
rect 3988 236132 3994 236134
rect 514017 232386 514083 232389
rect 583520 232386 584960 232476
rect 514017 232384 584960 232386
rect 514017 232328 514022 232384
rect 514078 232328 584960 232384
rect 514017 232326 584960 232328
rect 514017 232323 514083 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 514109 228034 514175 228037
rect 511796 228032 514175 228034
rect 511796 227976 514114 228032
rect 514170 227976 514175 228032
rect 511796 227974 514175 227976
rect 514109 227971 514175 227974
rect 580390 218996 580396 219060
rect 580460 219058 580466 219060
rect 583520 219058 584960 219148
rect 580460 218998 584960 219058
rect 580460 218996 580466 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 4061 214978 4127 214981
rect -960 214976 4127 214978
rect -960 214920 4066 214976
rect 4122 214920 4127 214976
rect -960 214918 4127 214920
rect -960 214828 480 214918
rect 4061 214915 4127 214918
rect 580206 205668 580212 205732
rect 580276 205730 580282 205732
rect 583520 205730 584960 205820
rect 580276 205670 584960 205730
rect 580276 205668 580282 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 514017 198114 514083 198117
rect 511796 198112 514083 198114
rect 511796 198056 514022 198112
rect 514078 198056 514083 198112
rect 511796 198054 514083 198056
rect 514017 198051 514083 198054
rect 514334 192476 514340 192540
rect 514404 192538 514410 192540
rect 583520 192538 584960 192628
rect 514404 192478 584960 192538
rect 514404 192476 514410 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 580206 179148 580212 179212
rect 580276 179210 580282 179212
rect 583520 179210 584960 179300
rect 580276 179150 584960 179210
rect 580276 179148 580282 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 3550 169492 3556 169556
rect 3620 169554 3626 169556
rect 3620 169494 12052 169554
rect 3620 169492 3626 169494
rect 580390 168194 580396 168196
rect 511796 168134 580396 168194
rect 580390 168132 580396 168134
rect 580460 168132 580466 168196
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 514201 152690 514267 152693
rect 583520 152690 584960 152780
rect 514201 152688 584960 152690
rect 514201 152632 514206 152688
rect 514262 152632 584960 152688
rect 514201 152630 584960 152632
rect 514201 152627 514267 152630
rect 583520 152540 584960 152630
rect -960 149684 480 149924
rect 580390 139300 580396 139364
rect 580460 139362 580466 139364
rect 583520 139362 584960 139452
rect 580460 139302 584960 139362
rect 580460 139300 580466 139302
rect 583520 139212 584960 139302
rect 580206 138274 580212 138276
rect 511796 138214 580212 138274
rect 580206 138212 580212 138214
rect 580276 138212 580282 138276
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 514150 112780 514156 112844
rect 514220 112842 514226 112844
rect 583520 112842 584960 112932
rect 514220 112782 584960 112842
rect 514220 112780 514226 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580390 108354 580396 108356
rect 511796 108294 580396 108354
rect 580390 108292 580396 108294
rect 580460 108292 580466 108356
rect 3734 102852 3740 102916
rect 3804 102914 3810 102916
rect 3804 102854 12052 102914
rect 3804 102852 3810 102854
rect 580206 99452 580212 99516
rect 580276 99514 580282 99516
rect 583520 99514 584960 99604
rect 580276 99454 584960 99514
rect 580276 99452 580282 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 580206 78434 580212 78436
rect 511796 78374 580212 78434
rect 580206 78372 580212 78374
rect 580276 78372 580282 78436
rect 514109 72994 514175 72997
rect 583520 72994 584960 73084
rect 514109 72992 584960 72994
rect 514109 72936 514114 72992
rect 514170 72936 584960 72992
rect 514109 72934 584960 72936
rect 514109 72931 514175 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2957 71634 3023 71637
rect -960 71632 3023 71634
rect -960 71576 2962 71632
rect 3018 71576 3023 71632
rect -960 71574 3023 71576
rect -960 71484 480 71574
rect 2957 71571 3023 71574
rect 580206 59604 580212 59668
rect 580276 59666 580282 59668
rect 583520 59666 584960 59756
rect 580276 59606 584960 59666
rect 580276 59604 580282 59606
rect 583520 59516 584960 59606
rect -960 58428 480 58668
rect 580206 48514 580212 48516
rect 511796 48454 580212 48514
rect 580206 48452 580212 48454
rect 580276 48452 580282 48516
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 3366 36212 3372 36276
rect 3436 36274 3442 36276
rect 3436 36214 12052 36274
rect 3436 36212 3442 36214
rect 514017 33146 514083 33149
rect 583520 33146 584960 33236
rect 514017 33144 584960 33146
rect 514017 33088 514022 33144
rect 514078 33088 584960 33144
rect 514017 33086 584960 33088
rect 514017 33083 514083 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 583520 19818 584960 19908
rect 518850 19758 584960 19818
rect -960 19260 480 19500
rect 518850 19410 518910 19758
rect 583520 19668 584960 19758
rect 513422 19350 518910 19410
rect 513422 19274 513482 19350
rect 511766 19214 513482 19274
rect 511766 18564 511826 19214
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 425375 3090 425441 3093
rect 580993 3090 581059 3093
rect 425375 3088 581059 3090
rect 425375 3032 425380 3088
rect 425436 3032 580998 3088
rect 581054 3032 581059 3088
rect 425375 3030 581059 3032
rect 425375 3027 425441 3030
rect 580993 3027 581059 3030
rect 463831 2954 463897 2957
rect 583385 2954 583451 2957
rect 463831 2952 583451 2954
rect 463831 2896 463836 2952
rect 463892 2896 583390 2952
rect 583446 2896 583451 2952
rect 463831 2894 583451 2896
rect 463831 2891 463897 2894
rect 583385 2891 583451 2894
rect 3141 1322 3207 1325
rect 252001 1322 252067 1325
rect 3141 1320 252067 1322
rect 3141 1264 3146 1320
rect 3202 1264 252006 1320
rect 252062 1264 252067 1320
rect 3141 1262 252067 1264
rect 3141 1259 3207 1262
rect 252001 1259 252067 1262
rect 271781 1322 271847 1325
rect 579797 1322 579863 1325
rect 271781 1320 579863 1322
rect 271781 1264 271786 1320
rect 271842 1264 579802 1320
rect 579858 1264 579863 1320
rect 271781 1262 579863 1264
rect 271781 1259 271847 1262
rect 579797 1259 579863 1262
rect 3325 1186 3391 1189
rect 232773 1186 232839 1189
rect 3325 1184 232839 1186
rect 3325 1128 3330 1184
rect 3386 1128 232778 1184
rect 232834 1128 232839 1184
rect 3325 1126 232839 1128
rect 3325 1123 3391 1126
rect 232773 1123 232839 1126
rect 291101 1186 291167 1189
rect 579981 1186 580047 1189
rect 291101 1184 580047 1186
rect 291101 1128 291106 1184
rect 291162 1128 579986 1184
rect 580042 1128 580047 1184
rect 291101 1126 580047 1128
rect 291101 1123 291167 1126
rect 579981 1123 580047 1126
rect 2957 1050 3023 1053
rect 59721 1050 59787 1053
rect 2957 1048 59787 1050
rect 2957 992 2962 1048
rect 3018 992 59726 1048
rect 59782 992 59787 1048
rect 2957 990 59787 992
rect 2957 987 3023 990
rect 59721 987 59787 990
rect 348785 1050 348851 1053
rect 580717 1050 580783 1053
rect 348785 1048 580783 1050
rect 348785 992 348790 1048
rect 348846 992 580722 1048
rect 580778 992 580783 1048
rect 348785 990 580783 992
rect 348785 987 348851 990
rect 580717 987 580783 990
rect 2773 914 2839 917
rect 40493 914 40559 917
rect 2773 912 40559 914
rect 2773 856 2778 912
rect 2834 856 40498 912
rect 40554 856 40559 912
rect 2773 854 40559 856
rect 2773 851 2839 854
rect 40493 851 40559 854
rect 98821 914 98887 917
rect 387701 914 387767 917
rect 98821 912 387767 914
rect 98821 856 98826 912
rect 98882 856 387706 912
rect 387762 856 387767 912
rect 98821 854 387767 856
rect 98821 851 98887 854
rect 387701 851 387767 854
rect 4061 778 4127 781
rect 213545 778 213611 781
rect 4061 776 213611 778
rect 4061 720 4066 776
rect 4122 720 213550 776
rect 213606 720 213611 776
rect 4061 718 213611 720
rect 4061 715 4127 718
rect 213545 715 213611 718
rect 310329 778 310395 781
rect 580165 778 580231 781
rect 310329 776 580231 778
rect 310329 720 310334 776
rect 310390 720 580170 776
rect 580226 720 580231 776
rect 310329 718 580231 720
rect 310329 715 310395 718
rect 580165 715 580231 718
rect 3877 642 3943 645
rect 194593 642 194659 645
rect 3877 640 194659 642
rect 3877 584 3882 640
rect 3938 584 194598 640
rect 194654 584 194659 640
rect 3877 582 194659 584
rect 3877 579 3943 582
rect 194593 579 194659 582
rect 329557 642 329623 645
rect 580901 642 580967 645
rect 329557 640 580967 642
rect 329557 584 329562 640
rect 329618 584 580906 640
rect 580962 584 580967 640
rect 329557 582 580967 584
rect 329557 579 329623 582
rect 580901 579 580967 582
rect 3693 506 3759 509
rect 175273 506 175339 509
rect 3693 504 175339 506
rect 3693 448 3698 504
rect 3754 448 175278 504
rect 175334 448 175339 504
rect 3693 446 175339 448
rect 3693 443 3759 446
rect 175273 443 175339 446
rect 368013 506 368079 509
rect 580533 506 580599 509
rect 368013 504 580599 506
rect 368013 448 368018 504
rect 368074 448 580538 504
rect 580594 448 580599 504
rect 368013 446 580599 448
rect 368013 443 368079 446
rect 580533 443 580599 446
rect 79501 370 79567 373
rect 368381 370 368447 373
rect 79501 368 368447 370
rect 79501 312 79506 368
rect 79562 312 368386 368
rect 368442 312 368447 368
rect 79501 310 368447 312
rect 79501 307 79567 310
rect 368381 307 368447 310
rect 386873 370 386939 373
rect 445661 370 445727 373
rect 386873 368 445727 370
rect 386873 312 386878 368
rect 386934 312 445666 368
rect 445722 312 445727 368
rect 386873 310 445727 312
rect 386873 307 386939 310
rect 445661 307 445727 310
rect 444833 98 444899 101
rect 581821 98 581887 101
rect 444833 96 581887 98
rect 444833 40 444838 96
rect 444894 40 581826 96
rect 581882 40 581887 96
rect 444833 38 581887 40
rect 444833 35 444899 38
rect 581821 35 581887 38
<< via3 >>
rect 3556 684252 3620 684316
rect 514156 643996 514220 644060
rect 3924 632028 3988 632092
rect 12020 602244 12084 602308
rect 580212 602244 580276 602308
rect 580396 590956 580460 591020
rect 514156 587012 514220 587076
rect 3372 579940 3436 580004
rect 12020 569332 12084 569396
rect 580396 557092 580460 557156
rect 514156 537780 514220 537844
rect 3740 527852 3804 527916
rect 514156 527172 514220 527236
rect 514156 497252 514220 497316
rect 514156 484604 514220 484668
rect 514340 467332 514404 467396
rect 514156 437412 514220 437476
rect 514340 431564 514404 431628
rect 514340 407492 514404 407556
rect 514156 378388 514220 378452
rect 514156 377572 514220 377636
rect 514340 325212 514404 325276
rect 514340 317732 514404 317796
rect 514156 272172 514220 272236
rect 514156 257892 514220 257956
rect 3924 236132 3988 236196
rect 580396 218996 580460 219060
rect 580212 205668 580276 205732
rect 514340 192476 514404 192540
rect 580212 179148 580276 179212
rect 3556 169492 3620 169556
rect 580396 168132 580460 168196
rect 580396 139300 580460 139364
rect 580212 138212 580276 138276
rect 514156 112780 514220 112844
rect 580396 108292 580460 108356
rect 3740 102852 3804 102916
rect 580212 99452 580276 99516
rect 580212 78372 580276 78436
rect 580212 59604 580276 59668
rect 580212 48452 580276 48516
rect 3372 36212 3436 36276
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3555 684316 3621 684317
rect 3555 684252 3556 684316
rect 3620 684252 3621 684316
rect 3555 684251 3621 684252
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3371 580004 3437 580005
rect 3371 579940 3372 580004
rect 3436 579940 3437 580004
rect 3371 579939 3437 579940
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 36277 3434 579939
rect 3558 169557 3618 684251
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 3923 632092 3989 632093
rect 3923 632028 3924 632092
rect 3988 632028 3989 632092
rect 3923 632027 3989 632028
rect 3739 527916 3805 527917
rect 3739 527852 3740 527916
rect 3804 527852 3805 527916
rect 3739 527851 3805 527852
rect 3555 169556 3621 169557
rect 3555 169492 3556 169556
rect 3620 169492 3621 169556
rect 3555 169491 3621 169492
rect 3742 102917 3802 527851
rect 3926 236197 3986 632027
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 3923 236196 3989 236197
rect 3923 236132 3924 236196
rect 3988 236132 3989 236196
rect 3923 236131 3989 236132
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3739 102916 3805 102917
rect 3739 102852 3740 102916
rect 3804 102852 3805 102916
rect 3739 102851 3805 102852
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 3371 36276 3437 36277
rect 3371 36212 3372 36276
rect 3436 36212 3437 36276
rect 3371 36211 3437 36212
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12019 602308 12085 602309
rect 12019 602244 12020 602308
rect 12084 602244 12085 602308
rect 12019 602243 12085 602244
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 12022 569397 12082 602243
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12019 569396 12085 569397
rect 12019 569332 12020 569396
rect 12084 569332 12085 569396
rect 12019 569331 12085 569332
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 554614 13574 590058
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16208 579454 16528 579486
rect 16208 579218 16250 579454
rect 16486 579218 16528 579454
rect 16208 579134 16528 579218
rect 16208 578898 16250 579134
rect 16486 578898 16528 579134
rect 16208 578866 16528 578898
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16208 543454 16528 543486
rect 16208 543218 16250 543454
rect 16486 543218 16528 543454
rect 16208 543134 16528 543218
rect 16208 542898 16250 543134
rect 16486 542898 16528 543134
rect 16208 542866 16528 542898
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16208 507454 16528 507486
rect 16208 507218 16250 507454
rect 16486 507218 16528 507454
rect 16208 507134 16528 507218
rect 16208 506898 16250 507134
rect 16486 506898 16528 507134
rect 16208 506866 16528 506898
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16208 471454 16528 471486
rect 16208 471218 16250 471454
rect 16486 471218 16528 471454
rect 16208 471134 16528 471218
rect 16208 470898 16250 471134
rect 16486 470898 16528 471134
rect 16208 470866 16528 470898
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16208 435454 16528 435486
rect 16208 435218 16250 435454
rect 16486 435218 16528 435454
rect 16208 435134 16528 435218
rect 16208 434898 16250 435134
rect 16486 434898 16528 435134
rect 16208 434866 16528 434898
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16208 399454 16528 399486
rect 16208 399218 16250 399454
rect 16486 399218 16528 399454
rect 16208 399134 16528 399218
rect 16208 398898 16250 399134
rect 16486 398898 16528 399134
rect 16208 398866 16528 398898
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16208 363454 16528 363486
rect 16208 363218 16250 363454
rect 16486 363218 16528 363454
rect 16208 363134 16528 363218
rect 16208 362898 16250 363134
rect 16486 362898 16528 363134
rect 16208 362866 16528 362898
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16208 327454 16528 327486
rect 16208 327218 16250 327454
rect 16486 327218 16528 327454
rect 16208 327134 16528 327218
rect 16208 326898 16250 327134
rect 16486 326898 16528 327134
rect 16208 326866 16528 326898
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16208 291454 16528 291486
rect 16208 291218 16250 291454
rect 16486 291218 16528 291454
rect 16208 291134 16528 291218
rect 16208 290898 16250 291134
rect 16486 290898 16528 291134
rect 16208 290866 16528 290898
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16208 255454 16528 255486
rect 16208 255218 16250 255454
rect 16486 255218 16528 255454
rect 16208 255134 16528 255218
rect 16208 254898 16250 255134
rect 16486 254898 16528 255134
rect 16208 254866 16528 254898
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16208 219454 16528 219486
rect 16208 219218 16250 219454
rect 16486 219218 16528 219454
rect 16208 219134 16528 219218
rect 16208 218898 16250 219134
rect 16486 218898 16528 219134
rect 16208 218866 16528 218898
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16208 183454 16528 183486
rect 16208 183218 16250 183454
rect 16486 183218 16528 183454
rect 16208 183134 16528 183218
rect 16208 182898 16250 183134
rect 16486 182898 16528 183134
rect 16208 182866 16528 182898
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16208 147454 16528 147486
rect 16208 147218 16250 147454
rect 16486 147218 16528 147454
rect 16208 147134 16528 147218
rect 16208 146898 16250 147134
rect 16486 146898 16528 147134
rect 16208 146866 16528 146898
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16208 111454 16528 111486
rect 16208 111218 16250 111454
rect 16486 111218 16528 111454
rect 16208 111134 16528 111218
rect 16208 110898 16250 111134
rect 16486 110898 16528 111134
rect 16208 110866 16528 110898
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16208 75454 16528 75486
rect 16208 75218 16250 75454
rect 16486 75218 16528 75454
rect 16208 75134 16528 75218
rect 16208 74898 16250 75134
rect 16486 74898 16528 75134
rect 16208 74866 16528 74898
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16208 39454 16528 39486
rect 16208 39218 16250 39454
rect 16486 39218 16528 39454
rect 16208 39134 16528 39218
rect 16208 38898 16250 39134
rect 16486 38898 16528 39134
rect 16208 38866 16528 38898
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 21328 583174 21648 583206
rect 21328 582938 21370 583174
rect 21606 582938 21648 583174
rect 21328 582854 21648 582938
rect 21328 582618 21370 582854
rect 21606 582618 21648 582854
rect 21328 582586 21648 582618
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 24114 565774 24734 601218
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 26448 586894 26768 586926
rect 26448 586658 26490 586894
rect 26726 586658 26768 586894
rect 26448 586574 26768 586658
rect 26448 586338 26490 586574
rect 26726 586338 26768 586574
rect 26448 586306 26768 586338
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 21328 547174 21648 547206
rect 21328 546938 21370 547174
rect 21606 546938 21648 547174
rect 21328 546854 21648 546938
rect 21328 546618 21370 546854
rect 21606 546618 21648 546854
rect 21328 546586 21648 546618
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 24114 529774 24734 565218
rect 27834 569494 28454 604938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 36688 594334 37008 594366
rect 36688 594098 36730 594334
rect 36966 594098 37008 594334
rect 36688 594014 37008 594098
rect 36688 593778 36730 594014
rect 36966 593778 37008 594014
rect 36688 593746 37008 593778
rect 31568 590614 31888 590646
rect 31568 590378 31610 590614
rect 31846 590378 31888 590614
rect 31568 590294 31888 590378
rect 31568 590058 31610 590294
rect 31846 590058 31888 590294
rect 31568 590026 31888 590058
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 26448 550894 26768 550926
rect 26448 550658 26490 550894
rect 26726 550658 26768 550894
rect 26448 550574 26768 550658
rect 26448 550338 26490 550574
rect 26726 550338 26768 550574
rect 26448 550306 26768 550338
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 21328 511174 21648 511206
rect 21328 510938 21370 511174
rect 21606 510938 21648 511174
rect 21328 510854 21648 510938
rect 21328 510618 21370 510854
rect 21606 510618 21648 510854
rect 21328 510586 21648 510618
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 24114 493774 24734 529218
rect 27834 533494 28454 568938
rect 37794 579454 38414 614898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 602500 42134 618618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 41808 598054 42128 598086
rect 41808 597818 41850 598054
rect 42086 597818 42128 598054
rect 41808 597734 42128 597818
rect 41808 597498 41850 597734
rect 42086 597498 42128 597734
rect 41808 597466 42128 597498
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 36688 558334 37008 558366
rect 36688 558098 36730 558334
rect 36966 558098 37008 558334
rect 36688 558014 37008 558098
rect 36688 557778 36730 558014
rect 36966 557778 37008 558014
rect 36688 557746 37008 557778
rect 31568 554614 31888 554646
rect 31568 554378 31610 554614
rect 31846 554378 31888 554614
rect 31568 554294 31888 554378
rect 31568 554058 31610 554294
rect 31846 554058 31888 554294
rect 31568 554026 31888 554058
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 26448 514894 26768 514926
rect 26448 514658 26490 514894
rect 26726 514658 26768 514894
rect 26448 514574 26768 514658
rect 26448 514338 26490 514574
rect 26726 514338 26768 514574
rect 26448 514306 26768 514338
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 21328 475174 21648 475206
rect 21328 474938 21370 475174
rect 21606 474938 21648 475174
rect 21328 474854 21648 474938
rect 21328 474618 21370 474854
rect 21606 474618 21648 474854
rect 21328 474586 21648 474618
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 24114 457774 24734 493218
rect 27834 497494 28454 532938
rect 37794 543454 38414 578898
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 41808 562054 42128 562086
rect 41808 561818 41850 562054
rect 42086 561818 42128 562054
rect 41808 561734 42128 561818
rect 41808 561498 41850 561734
rect 42086 561498 42128 561734
rect 41808 561466 42128 561498
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 36688 522334 37008 522366
rect 36688 522098 36730 522334
rect 36966 522098 37008 522334
rect 36688 522014 37008 522098
rect 36688 521778 36730 522014
rect 36966 521778 37008 522014
rect 36688 521746 37008 521778
rect 31568 518614 31888 518646
rect 31568 518378 31610 518614
rect 31846 518378 31888 518614
rect 31568 518294 31888 518378
rect 31568 518058 31610 518294
rect 31846 518058 31888 518294
rect 31568 518026 31888 518058
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 26448 478894 26768 478926
rect 26448 478658 26490 478894
rect 26726 478658 26768 478894
rect 26448 478574 26768 478658
rect 26448 478338 26490 478574
rect 26726 478338 26768 478574
rect 26448 478306 26768 478338
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 21328 439174 21648 439206
rect 21328 438938 21370 439174
rect 21606 438938 21648 439174
rect 21328 438854 21648 438938
rect 21328 438618 21370 438854
rect 21606 438618 21648 438854
rect 21328 438586 21648 438618
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 24114 421774 24734 457218
rect 27834 461494 28454 496938
rect 37794 507454 38414 542898
rect 45234 550894 45854 586338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 46928 579454 47248 579486
rect 46928 579218 46970 579454
rect 47206 579218 47248 579454
rect 46928 579134 47248 579218
rect 46928 578898 46970 579134
rect 47206 578898 47248 579134
rect 46928 578866 47248 578898
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 41808 526054 42128 526086
rect 41808 525818 41850 526054
rect 42086 525818 42128 526054
rect 41808 525734 42128 525818
rect 41808 525498 41850 525734
rect 42086 525498 42128 525734
rect 41808 525466 42128 525498
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 36688 486334 37008 486366
rect 36688 486098 36730 486334
rect 36966 486098 37008 486334
rect 36688 486014 37008 486098
rect 36688 485778 36730 486014
rect 36966 485778 37008 486014
rect 36688 485746 37008 485778
rect 31568 482614 31888 482646
rect 31568 482378 31610 482614
rect 31846 482378 31888 482614
rect 31568 482294 31888 482378
rect 31568 482058 31610 482294
rect 31846 482058 31888 482294
rect 31568 482026 31888 482058
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 26448 442894 26768 442926
rect 26448 442658 26490 442894
rect 26726 442658 26768 442894
rect 26448 442574 26768 442658
rect 26448 442338 26490 442574
rect 26726 442338 26768 442574
rect 26448 442306 26768 442338
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 21328 403174 21648 403206
rect 21328 402938 21370 403174
rect 21606 402938 21648 403174
rect 21328 402854 21648 402938
rect 21328 402618 21370 402854
rect 21606 402618 21648 402854
rect 21328 402586 21648 402618
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 24114 385774 24734 421218
rect 27834 425494 28454 460938
rect 37794 471454 38414 506898
rect 45234 514894 45854 550338
rect 48954 554614 49574 590058
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52048 583174 52368 583206
rect 52048 582938 52090 583174
rect 52326 582938 52368 583174
rect 52048 582854 52368 582938
rect 52048 582618 52090 582854
rect 52326 582618 52368 582854
rect 52048 582586 52368 582618
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 46928 543454 47248 543486
rect 46928 543218 46970 543454
rect 47206 543218 47248 543454
rect 46928 543134 47248 543218
rect 46928 542898 46970 543134
rect 47206 542898 47248 543134
rect 46928 542866 47248 542898
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 41808 490054 42128 490086
rect 41808 489818 41850 490054
rect 42086 489818 42128 490054
rect 41808 489734 42128 489818
rect 41808 489498 41850 489734
rect 42086 489498 42128 489734
rect 41808 489466 42128 489498
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 36688 450334 37008 450366
rect 36688 450098 36730 450334
rect 36966 450098 37008 450334
rect 36688 450014 37008 450098
rect 36688 449778 36730 450014
rect 36966 449778 37008 450014
rect 36688 449746 37008 449778
rect 31568 446614 31888 446646
rect 31568 446378 31610 446614
rect 31846 446378 31888 446614
rect 31568 446294 31888 446378
rect 31568 446058 31610 446294
rect 31846 446058 31888 446294
rect 31568 446026 31888 446058
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 26448 406894 26768 406926
rect 26448 406658 26490 406894
rect 26726 406658 26768 406894
rect 26448 406574 26768 406658
rect 26448 406338 26490 406574
rect 26726 406338 26768 406574
rect 26448 406306 26768 406338
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 21328 367174 21648 367206
rect 21328 366938 21370 367174
rect 21606 366938 21648 367174
rect 21328 366854 21648 366938
rect 21328 366618 21370 366854
rect 21606 366618 21648 366854
rect 21328 366586 21648 366618
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 24114 349774 24734 385218
rect 27834 389494 28454 424938
rect 37794 435454 38414 470898
rect 45234 478894 45854 514338
rect 48954 518614 49574 554058
rect 52674 558334 53294 593778
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52048 547174 52368 547206
rect 52048 546938 52090 547174
rect 52326 546938 52368 547174
rect 52048 546854 52368 546938
rect 52048 546618 52090 546854
rect 52326 546618 52368 546854
rect 52048 546586 52368 546618
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 46928 507454 47248 507486
rect 46928 507218 46970 507454
rect 47206 507218 47248 507454
rect 46928 507134 47248 507218
rect 46928 506898 46970 507134
rect 47206 506898 47248 507134
rect 46928 506866 47248 506898
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 41808 454054 42128 454086
rect 41808 453818 41850 454054
rect 42086 453818 42128 454054
rect 41808 453734 42128 453818
rect 41808 453498 41850 453734
rect 42086 453498 42128 453734
rect 41808 453466 42128 453498
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 36688 414334 37008 414366
rect 36688 414098 36730 414334
rect 36966 414098 37008 414334
rect 36688 414014 37008 414098
rect 36688 413778 36730 414014
rect 36966 413778 37008 414014
rect 36688 413746 37008 413778
rect 31568 410614 31888 410646
rect 31568 410378 31610 410614
rect 31846 410378 31888 410614
rect 31568 410294 31888 410378
rect 31568 410058 31610 410294
rect 31846 410058 31888 410294
rect 31568 410026 31888 410058
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 26448 370894 26768 370926
rect 26448 370658 26490 370894
rect 26726 370658 26768 370894
rect 26448 370574 26768 370658
rect 26448 370338 26490 370574
rect 26726 370338 26768 370574
rect 26448 370306 26768 370338
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 21328 331174 21648 331206
rect 21328 330938 21370 331174
rect 21606 330938 21648 331174
rect 21328 330854 21648 330938
rect 21328 330618 21370 330854
rect 21606 330618 21648 330854
rect 21328 330586 21648 330618
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 24114 313774 24734 349218
rect 27834 353494 28454 388938
rect 37794 399454 38414 434898
rect 45234 442894 45854 478338
rect 48954 482614 49574 518058
rect 52674 522334 53294 557778
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52048 511174 52368 511206
rect 52048 510938 52090 511174
rect 52326 510938 52368 511174
rect 52048 510854 52368 510938
rect 52048 510618 52090 510854
rect 52326 510618 52368 510854
rect 52048 510586 52368 510618
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 46928 471454 47248 471486
rect 46928 471218 46970 471454
rect 47206 471218 47248 471454
rect 46928 471134 47248 471218
rect 46928 470898 46970 471134
rect 47206 470898 47248 471134
rect 46928 470866 47248 470898
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 41808 418054 42128 418086
rect 41808 417818 41850 418054
rect 42086 417818 42128 418054
rect 41808 417734 42128 417818
rect 41808 417498 41850 417734
rect 42086 417498 42128 417734
rect 41808 417466 42128 417498
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 36688 378334 37008 378366
rect 36688 378098 36730 378334
rect 36966 378098 37008 378334
rect 36688 378014 37008 378098
rect 36688 377778 36730 378014
rect 36966 377778 37008 378014
rect 36688 377746 37008 377778
rect 31568 374614 31888 374646
rect 31568 374378 31610 374614
rect 31846 374378 31888 374614
rect 31568 374294 31888 374378
rect 31568 374058 31610 374294
rect 31846 374058 31888 374294
rect 31568 374026 31888 374058
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 26448 334894 26768 334926
rect 26448 334658 26490 334894
rect 26726 334658 26768 334894
rect 26448 334574 26768 334658
rect 26448 334338 26490 334574
rect 26726 334338 26768 334574
rect 26448 334306 26768 334338
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 21328 295174 21648 295206
rect 21328 294938 21370 295174
rect 21606 294938 21648 295174
rect 21328 294854 21648 294938
rect 21328 294618 21370 294854
rect 21606 294618 21648 294854
rect 21328 294586 21648 294618
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 24114 277774 24734 313218
rect 27834 317494 28454 352938
rect 37794 363454 38414 398898
rect 45234 406894 45854 442338
rect 48954 446614 49574 482058
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52048 475174 52368 475206
rect 52048 474938 52090 475174
rect 52326 474938 52368 475174
rect 52048 474854 52368 474938
rect 52048 474618 52090 474854
rect 52326 474618 52368 474854
rect 52048 474586 52368 474618
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 46928 435454 47248 435486
rect 46928 435218 46970 435454
rect 47206 435218 47248 435454
rect 46928 435134 47248 435218
rect 46928 434898 46970 435134
rect 47206 434898 47248 435134
rect 46928 434866 47248 434898
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 41808 382054 42128 382086
rect 41808 381818 41850 382054
rect 42086 381818 42128 382054
rect 41808 381734 42128 381818
rect 41808 381498 41850 381734
rect 42086 381498 42128 381734
rect 41808 381466 42128 381498
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 36688 342334 37008 342366
rect 36688 342098 36730 342334
rect 36966 342098 37008 342334
rect 36688 342014 37008 342098
rect 36688 341778 36730 342014
rect 36966 341778 37008 342014
rect 36688 341746 37008 341778
rect 31568 338614 31888 338646
rect 31568 338378 31610 338614
rect 31846 338378 31888 338614
rect 31568 338294 31888 338378
rect 31568 338058 31610 338294
rect 31846 338058 31888 338294
rect 31568 338026 31888 338058
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 26448 298894 26768 298926
rect 26448 298658 26490 298894
rect 26726 298658 26768 298894
rect 26448 298574 26768 298658
rect 26448 298338 26490 298574
rect 26726 298338 26768 298574
rect 26448 298306 26768 298338
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 21328 259174 21648 259206
rect 21328 258938 21370 259174
rect 21606 258938 21648 259174
rect 21328 258854 21648 258938
rect 21328 258618 21370 258854
rect 21606 258618 21648 258854
rect 21328 258586 21648 258618
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 24114 241774 24734 277218
rect 27834 281494 28454 316938
rect 37794 327454 38414 362898
rect 45234 370894 45854 406338
rect 48954 410614 49574 446058
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52048 439174 52368 439206
rect 52048 438938 52090 439174
rect 52326 438938 52368 439174
rect 52048 438854 52368 438938
rect 52048 438618 52090 438854
rect 52326 438618 52368 438854
rect 52048 438586 52368 438618
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 46928 399454 47248 399486
rect 46928 399218 46970 399454
rect 47206 399218 47248 399454
rect 46928 399134 47248 399218
rect 46928 398898 46970 399134
rect 47206 398898 47248 399134
rect 46928 398866 47248 398898
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 41808 346054 42128 346086
rect 41808 345818 41850 346054
rect 42086 345818 42128 346054
rect 41808 345734 42128 345818
rect 41808 345498 41850 345734
rect 42086 345498 42128 345734
rect 41808 345466 42128 345498
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 36688 306334 37008 306366
rect 36688 306098 36730 306334
rect 36966 306098 37008 306334
rect 36688 306014 37008 306098
rect 36688 305778 36730 306014
rect 36966 305778 37008 306014
rect 36688 305746 37008 305778
rect 31568 302614 31888 302646
rect 31568 302378 31610 302614
rect 31846 302378 31888 302614
rect 31568 302294 31888 302378
rect 31568 302058 31610 302294
rect 31846 302058 31888 302294
rect 31568 302026 31888 302058
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 26448 262894 26768 262926
rect 26448 262658 26490 262894
rect 26726 262658 26768 262894
rect 26448 262574 26768 262658
rect 26448 262338 26490 262574
rect 26726 262338 26768 262574
rect 26448 262306 26768 262338
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 21328 223174 21648 223206
rect 21328 222938 21370 223174
rect 21606 222938 21648 223174
rect 21328 222854 21648 222938
rect 21328 222618 21370 222854
rect 21606 222618 21648 222854
rect 21328 222586 21648 222618
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 24114 205774 24734 241218
rect 27834 245494 28454 280938
rect 37794 291454 38414 326898
rect 45234 334894 45854 370338
rect 48954 374614 49574 410058
rect 52674 414334 53294 449778
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52048 403174 52368 403206
rect 52048 402938 52090 403174
rect 52326 402938 52368 403174
rect 52048 402854 52368 402938
rect 52048 402618 52090 402854
rect 52326 402618 52368 402854
rect 52048 402586 52368 402618
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 46928 363454 47248 363486
rect 46928 363218 46970 363454
rect 47206 363218 47248 363454
rect 46928 363134 47248 363218
rect 46928 362898 46970 363134
rect 47206 362898 47248 363134
rect 46928 362866 47248 362898
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 41808 310054 42128 310086
rect 41808 309818 41850 310054
rect 42086 309818 42128 310054
rect 41808 309734 42128 309818
rect 41808 309498 41850 309734
rect 42086 309498 42128 309734
rect 41808 309466 42128 309498
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 36688 270334 37008 270366
rect 36688 270098 36730 270334
rect 36966 270098 37008 270334
rect 36688 270014 37008 270098
rect 36688 269778 36730 270014
rect 36966 269778 37008 270014
rect 36688 269746 37008 269778
rect 31568 266614 31888 266646
rect 31568 266378 31610 266614
rect 31846 266378 31888 266614
rect 31568 266294 31888 266378
rect 31568 266058 31610 266294
rect 31846 266058 31888 266294
rect 31568 266026 31888 266058
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 26448 226894 26768 226926
rect 26448 226658 26490 226894
rect 26726 226658 26768 226894
rect 26448 226574 26768 226658
rect 26448 226338 26490 226574
rect 26726 226338 26768 226574
rect 26448 226306 26768 226338
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 21328 187174 21648 187206
rect 21328 186938 21370 187174
rect 21606 186938 21648 187174
rect 21328 186854 21648 186938
rect 21328 186618 21370 186854
rect 21606 186618 21648 186854
rect 21328 186586 21648 186618
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 24114 169774 24734 205218
rect 27834 209494 28454 244938
rect 37794 255454 38414 290898
rect 45234 298894 45854 334338
rect 48954 338614 49574 374058
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52048 367174 52368 367206
rect 52048 366938 52090 367174
rect 52326 366938 52368 367174
rect 52048 366854 52368 366938
rect 52048 366618 52090 366854
rect 52326 366618 52368 366854
rect 52048 366586 52368 366618
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 46928 327454 47248 327486
rect 46928 327218 46970 327454
rect 47206 327218 47248 327454
rect 46928 327134 47248 327218
rect 46928 326898 46970 327134
rect 47206 326898 47248 327134
rect 46928 326866 47248 326898
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 41808 274054 42128 274086
rect 41808 273818 41850 274054
rect 42086 273818 42128 274054
rect 41808 273734 42128 273818
rect 41808 273498 41850 273734
rect 42086 273498 42128 273734
rect 41808 273466 42128 273498
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 36688 234334 37008 234366
rect 36688 234098 36730 234334
rect 36966 234098 37008 234334
rect 36688 234014 37008 234098
rect 36688 233778 36730 234014
rect 36966 233778 37008 234014
rect 36688 233746 37008 233778
rect 31568 230614 31888 230646
rect 31568 230378 31610 230614
rect 31846 230378 31888 230614
rect 31568 230294 31888 230378
rect 31568 230058 31610 230294
rect 31846 230058 31888 230294
rect 31568 230026 31888 230058
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 26448 190894 26768 190926
rect 26448 190658 26490 190894
rect 26726 190658 26768 190894
rect 26448 190574 26768 190658
rect 26448 190338 26490 190574
rect 26726 190338 26768 190574
rect 26448 190306 26768 190338
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 21328 151174 21648 151206
rect 21328 150938 21370 151174
rect 21606 150938 21648 151174
rect 21328 150854 21648 150938
rect 21328 150618 21370 150854
rect 21606 150618 21648 150854
rect 21328 150586 21648 150618
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 24114 133774 24734 169218
rect 27834 173494 28454 208938
rect 37794 219454 38414 254898
rect 45234 262894 45854 298338
rect 48954 302614 49574 338058
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52048 331174 52368 331206
rect 52048 330938 52090 331174
rect 52326 330938 52368 331174
rect 52048 330854 52368 330938
rect 52048 330618 52090 330854
rect 52326 330618 52368 330854
rect 52048 330586 52368 330618
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 46928 291454 47248 291486
rect 46928 291218 46970 291454
rect 47206 291218 47248 291454
rect 46928 291134 47248 291218
rect 46928 290898 46970 291134
rect 47206 290898 47248 291134
rect 46928 290866 47248 290898
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 41808 238054 42128 238086
rect 41808 237818 41850 238054
rect 42086 237818 42128 238054
rect 41808 237734 42128 237818
rect 41808 237498 41850 237734
rect 42086 237498 42128 237734
rect 41808 237466 42128 237498
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 36688 198334 37008 198366
rect 36688 198098 36730 198334
rect 36966 198098 37008 198334
rect 36688 198014 37008 198098
rect 36688 197778 36730 198014
rect 36966 197778 37008 198014
rect 36688 197746 37008 197778
rect 31568 194614 31888 194646
rect 31568 194378 31610 194614
rect 31846 194378 31888 194614
rect 31568 194294 31888 194378
rect 31568 194058 31610 194294
rect 31846 194058 31888 194294
rect 31568 194026 31888 194058
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 26448 154894 26768 154926
rect 26448 154658 26490 154894
rect 26726 154658 26768 154894
rect 26448 154574 26768 154658
rect 26448 154338 26490 154574
rect 26726 154338 26768 154574
rect 26448 154306 26768 154338
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 21328 115174 21648 115206
rect 21328 114938 21370 115174
rect 21606 114938 21648 115174
rect 21328 114854 21648 114938
rect 21328 114618 21370 114854
rect 21606 114618 21648 114854
rect 21328 114586 21648 114618
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 24114 97774 24734 133218
rect 27834 137494 28454 172938
rect 37794 183454 38414 218898
rect 45234 226894 45854 262338
rect 48954 266614 49574 302058
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52048 295174 52368 295206
rect 52048 294938 52090 295174
rect 52326 294938 52368 295174
rect 52048 294854 52368 294938
rect 52048 294618 52090 294854
rect 52326 294618 52368 294854
rect 52048 294586 52368 294618
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 46928 255454 47248 255486
rect 46928 255218 46970 255454
rect 47206 255218 47248 255454
rect 46928 255134 47248 255218
rect 46928 254898 46970 255134
rect 47206 254898 47248 255134
rect 46928 254866 47248 254898
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 41808 202054 42128 202086
rect 41808 201818 41850 202054
rect 42086 201818 42128 202054
rect 41808 201734 42128 201818
rect 41808 201498 41850 201734
rect 42086 201498 42128 201734
rect 41808 201466 42128 201498
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 36688 162334 37008 162366
rect 36688 162098 36730 162334
rect 36966 162098 37008 162334
rect 36688 162014 37008 162098
rect 36688 161778 36730 162014
rect 36966 161778 37008 162014
rect 36688 161746 37008 161778
rect 31568 158614 31888 158646
rect 31568 158378 31610 158614
rect 31846 158378 31888 158614
rect 31568 158294 31888 158378
rect 31568 158058 31610 158294
rect 31846 158058 31888 158294
rect 31568 158026 31888 158058
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 26448 118894 26768 118926
rect 26448 118658 26490 118894
rect 26726 118658 26768 118894
rect 26448 118574 26768 118658
rect 26448 118338 26490 118574
rect 26726 118338 26768 118574
rect 26448 118306 26768 118338
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 21328 79174 21648 79206
rect 21328 78938 21370 79174
rect 21606 78938 21648 79174
rect 21328 78854 21648 78938
rect 21328 78618 21370 78854
rect 21606 78618 21648 78854
rect 21328 78586 21648 78618
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 24114 61774 24734 97218
rect 27834 101494 28454 136938
rect 37794 147454 38414 182898
rect 45234 190894 45854 226338
rect 48954 230614 49574 266058
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52048 259174 52368 259206
rect 52048 258938 52090 259174
rect 52326 258938 52368 259174
rect 52048 258854 52368 258938
rect 52048 258618 52090 258854
rect 52326 258618 52368 258854
rect 52048 258586 52368 258618
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 46928 219454 47248 219486
rect 46928 219218 46970 219454
rect 47206 219218 47248 219454
rect 46928 219134 47248 219218
rect 46928 218898 46970 219134
rect 47206 218898 47248 219134
rect 46928 218866 47248 218898
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 41808 166054 42128 166086
rect 41808 165818 41850 166054
rect 42086 165818 42128 166054
rect 41808 165734 42128 165818
rect 41808 165498 41850 165734
rect 42086 165498 42128 165734
rect 41808 165466 42128 165498
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 36688 126334 37008 126366
rect 36688 126098 36730 126334
rect 36966 126098 37008 126334
rect 36688 126014 37008 126098
rect 36688 125778 36730 126014
rect 36966 125778 37008 126014
rect 36688 125746 37008 125778
rect 31568 122614 31888 122646
rect 31568 122378 31610 122614
rect 31846 122378 31888 122614
rect 31568 122294 31888 122378
rect 31568 122058 31610 122294
rect 31846 122058 31888 122294
rect 31568 122026 31888 122058
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 26448 82894 26768 82926
rect 26448 82658 26490 82894
rect 26726 82658 26768 82894
rect 26448 82574 26768 82658
rect 26448 82338 26490 82574
rect 26726 82338 26768 82574
rect 26448 82306 26768 82338
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 21328 43174 21648 43206
rect 21328 42938 21370 43174
rect 21606 42938 21648 43174
rect 21328 42854 21648 42938
rect 21328 42618 21370 42854
rect 21606 42618 21648 42854
rect 21328 42586 21648 42618
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 24114 25774 24734 61218
rect 27834 65494 28454 100938
rect 37794 111454 38414 146898
rect 45234 154894 45854 190338
rect 48954 194614 49574 230058
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52048 223174 52368 223206
rect 52048 222938 52090 223174
rect 52326 222938 52368 223174
rect 52048 222854 52368 222938
rect 52048 222618 52090 222854
rect 52326 222618 52368 222854
rect 52048 222586 52368 222618
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 46928 183454 47248 183486
rect 46928 183218 46970 183454
rect 47206 183218 47248 183454
rect 46928 183134 47248 183218
rect 46928 182898 46970 183134
rect 47206 182898 47248 183134
rect 46928 182866 47248 182898
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 41808 130054 42128 130086
rect 41808 129818 41850 130054
rect 42086 129818 42128 130054
rect 41808 129734 42128 129818
rect 41808 129498 41850 129734
rect 42086 129498 42128 129734
rect 41808 129466 42128 129498
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 36688 90334 37008 90366
rect 36688 90098 36730 90334
rect 36966 90098 37008 90334
rect 36688 90014 37008 90098
rect 36688 89778 36730 90014
rect 36966 89778 37008 90014
rect 36688 89746 37008 89778
rect 31568 86614 31888 86646
rect 31568 86378 31610 86614
rect 31846 86378 31888 86614
rect 31568 86294 31888 86378
rect 31568 86058 31610 86294
rect 31846 86058 31888 86294
rect 31568 86026 31888 86058
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 26448 46894 26768 46926
rect 26448 46658 26490 46894
rect 26726 46658 26768 46894
rect 26448 46574 26768 46658
rect 26448 46338 26490 46574
rect 26726 46338 26768 46574
rect 26448 46306 26768 46338
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 21328 7174 21648 7206
rect 21328 6938 21370 7174
rect 21606 6938 21648 7174
rect 21328 6854 21648 6938
rect 21328 6618 21370 6854
rect 21606 6618 21648 6854
rect 21328 6586 21648 6618
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 -6106 24734 25218
rect 27834 29494 28454 64938
rect 37794 75454 38414 110898
rect 45234 118894 45854 154338
rect 48954 158614 49574 194058
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52048 187174 52368 187206
rect 52048 186938 52090 187174
rect 52326 186938 52368 187174
rect 52048 186854 52368 186938
rect 52048 186618 52090 186854
rect 52326 186618 52368 186854
rect 52048 186586 52368 186618
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 46928 147454 47248 147486
rect 46928 147218 46970 147454
rect 47206 147218 47248 147454
rect 46928 147134 47248 147218
rect 46928 146898 46970 147134
rect 47206 146898 47248 147134
rect 46928 146866 47248 146898
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 41808 94054 42128 94086
rect 41808 93818 41850 94054
rect 42086 93818 42128 94054
rect 41808 93734 42128 93818
rect 41808 93498 41850 93734
rect 42086 93498 42128 93734
rect 41808 93466 42128 93498
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 36688 54334 37008 54366
rect 36688 54098 36730 54334
rect 36966 54098 37008 54334
rect 36688 54014 37008 54098
rect 36688 53778 36730 54014
rect 36966 53778 37008 54014
rect 36688 53746 37008 53778
rect 31568 50614 31888 50646
rect 31568 50378 31610 50614
rect 31846 50378 31888 50614
rect 31568 50294 31888 50378
rect 31568 50058 31610 50294
rect 31846 50058 31888 50294
rect 31568 50026 31888 50058
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 26448 10894 26768 10926
rect 26448 10658 26490 10894
rect 26726 10658 26768 10894
rect 26448 10574 26768 10658
rect 26448 10338 26490 10574
rect 26726 10338 26768 10574
rect 26448 10306 26768 10338
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 -7066 28454 28938
rect 37794 39454 38414 74898
rect 45234 82894 45854 118338
rect 48954 122614 49574 158058
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52048 151174 52368 151206
rect 52048 150938 52090 151174
rect 52326 150938 52368 151174
rect 52048 150854 52368 150938
rect 52048 150618 52090 150854
rect 52326 150618 52368 150854
rect 52048 150586 52368 150618
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 46928 111454 47248 111486
rect 46928 111218 46970 111454
rect 47206 111218 47248 111454
rect 46928 111134 47248 111218
rect 46928 110898 46970 111134
rect 47206 110898 47248 111134
rect 46928 110866 47248 110898
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 41808 58054 42128 58086
rect 41808 57818 41850 58054
rect 42086 57818 42128 58054
rect 41808 57734 42128 57818
rect 41808 57498 41850 57734
rect 42086 57498 42128 57734
rect 41808 57466 42128 57498
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 36688 18334 37008 18366
rect 36688 18098 36730 18334
rect 36966 18098 37008 18334
rect 36688 18014 37008 18098
rect 36688 17778 36730 18014
rect 36966 17778 37008 18014
rect 36688 17746 37008 17778
rect 31568 14614 31888 14646
rect 31568 14378 31610 14614
rect 31846 14378 31888 14614
rect 31568 14294 31888 14378
rect 31568 14058 31610 14294
rect 31846 14058 31888 14294
rect 31568 14026 31888 14058
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 3454 38414 38898
rect 45234 46894 45854 82338
rect 48954 86614 49574 122058
rect 52674 126334 53294 161778
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52048 115174 52368 115206
rect 52048 114938 52090 115174
rect 52326 114938 52368 115174
rect 52048 114854 52368 114938
rect 52048 114618 52090 114854
rect 52326 114618 52368 114854
rect 52048 114586 52368 114618
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 46928 75454 47248 75486
rect 46928 75218 46970 75454
rect 47206 75218 47248 75454
rect 46928 75134 47248 75218
rect 46928 74898 46970 75134
rect 47206 74898 47248 75134
rect 46928 74866 47248 74898
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 41808 22054 42128 22086
rect 41808 21818 41850 22054
rect 42086 21818 42128 22054
rect 41808 21734 42128 21818
rect 41808 21498 41850 21734
rect 42086 21498 42128 21734
rect 41808 21466 42128 21498
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 45234 10894 45854 46338
rect 48954 50614 49574 86058
rect 52674 90334 53294 125778
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52048 79174 52368 79206
rect 52048 78938 52090 79174
rect 52326 78938 52368 79174
rect 52048 78854 52368 78938
rect 52048 78618 52090 78854
rect 52326 78618 52368 78854
rect 52048 78586 52368 78618
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 46928 39454 47248 39486
rect 46928 39218 46970 39454
rect 47206 39218 47248 39454
rect 46928 39134 47248 39218
rect 46928 38898 46970 39134
rect 47206 38898 47248 39134
rect 46928 38866 47248 38898
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 -1306 42134 2988
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 50058
rect 52674 54334 53294 89778
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52048 43174 52368 43206
rect 52048 42938 52090 43174
rect 52326 42938 52368 43174
rect 52048 42854 52368 42938
rect 52048 42618 52090 42854
rect 52326 42618 52368 42854
rect 52048 42586 52368 42618
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52048 7174 52368 7206
rect 52048 6938 52090 7174
rect 52326 6938 52368 7174
rect 52048 6854 52368 6938
rect 52048 6618 52090 6854
rect 52326 6618 52368 6854
rect 52048 6586 52368 6618
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 57168 586894 57488 586926
rect 57168 586658 57210 586894
rect 57446 586658 57488 586894
rect 57168 586574 57488 586658
rect 57168 586338 57210 586574
rect 57446 586338 57488 586574
rect 57168 586306 57488 586338
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 56394 526054 57014 561498
rect 60114 565774 60734 601218
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 605494 64454 640938
rect 63834 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 64454 605494
rect 63834 605174 64454 605258
rect 63834 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 64454 605174
rect 62288 590614 62608 590646
rect 62288 590378 62330 590614
rect 62566 590378 62608 590614
rect 62288 590294 62608 590378
rect 62288 590058 62330 590294
rect 62566 590058 62608 590294
rect 62288 590026 62608 590058
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 57168 550894 57488 550926
rect 57168 550658 57210 550894
rect 57446 550658 57488 550894
rect 57168 550574 57488 550658
rect 57168 550338 57210 550574
rect 57446 550338 57488 550574
rect 57168 550306 57488 550338
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 56394 490054 57014 525498
rect 60114 529774 60734 565218
rect 63834 569494 64454 604938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 72528 598054 72848 598086
rect 72528 597818 72570 598054
rect 72806 597818 72848 598054
rect 72528 597734 72848 597818
rect 72528 597498 72570 597734
rect 72806 597498 72848 597734
rect 72528 597466 72848 597498
rect 67408 594334 67728 594366
rect 67408 594098 67450 594334
rect 67686 594098 67728 594334
rect 67408 594014 67728 594098
rect 67408 593778 67450 594014
rect 67686 593778 67728 594014
rect 67408 593746 67728 593778
rect 63834 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 64454 569494
rect 63834 569174 64454 569258
rect 63834 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 64454 569174
rect 62288 554614 62608 554646
rect 62288 554378 62330 554614
rect 62566 554378 62608 554614
rect 62288 554294 62608 554378
rect 62288 554058 62330 554294
rect 62566 554058 62608 554294
rect 62288 554026 62608 554058
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 57168 514894 57488 514926
rect 57168 514658 57210 514894
rect 57446 514658 57488 514894
rect 57168 514574 57488 514658
rect 57168 514338 57210 514574
rect 57446 514338 57488 514574
rect 57168 514306 57488 514338
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 60114 493774 60734 529218
rect 63834 533494 64454 568938
rect 73794 579454 74414 614898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 602500 78134 618618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 72528 562054 72848 562086
rect 72528 561818 72570 562054
rect 72806 561818 72848 562054
rect 72528 561734 72848 561818
rect 72528 561498 72570 561734
rect 72806 561498 72848 561734
rect 72528 561466 72848 561498
rect 67408 558334 67728 558366
rect 67408 558098 67450 558334
rect 67686 558098 67728 558334
rect 67408 558014 67728 558098
rect 67408 557778 67450 558014
rect 67686 557778 67728 558014
rect 67408 557746 67728 557778
rect 63834 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 64454 533494
rect 63834 533174 64454 533258
rect 63834 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 64454 533174
rect 62288 518614 62608 518646
rect 62288 518378 62330 518614
rect 62566 518378 62608 518614
rect 62288 518294 62608 518378
rect 62288 518058 62330 518294
rect 62566 518058 62608 518294
rect 62288 518026 62608 518058
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 57168 478894 57488 478926
rect 57168 478658 57210 478894
rect 57446 478658 57488 478894
rect 57168 478574 57488 478658
rect 57168 478338 57210 478574
rect 57446 478338 57488 478574
rect 57168 478306 57488 478338
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 60114 457774 60734 493218
rect 63834 497494 64454 532938
rect 73794 543454 74414 578898
rect 77648 579454 77968 579486
rect 77648 579218 77690 579454
rect 77926 579218 77968 579454
rect 77648 579134 77968 579218
rect 77648 578898 77690 579134
rect 77926 578898 77968 579134
rect 77648 578866 77968 578898
rect 81234 550894 81854 586338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 82768 583174 83088 583206
rect 82768 582938 82810 583174
rect 83046 582938 83088 583174
rect 82768 582854 83088 582938
rect 82768 582618 82810 582854
rect 83046 582618 83088 582854
rect 82768 582586 83088 582618
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 72528 526054 72848 526086
rect 72528 525818 72570 526054
rect 72806 525818 72848 526054
rect 72528 525734 72848 525818
rect 72528 525498 72570 525734
rect 72806 525498 72848 525734
rect 72528 525466 72848 525498
rect 67408 522334 67728 522366
rect 67408 522098 67450 522334
rect 67686 522098 67728 522334
rect 67408 522014 67728 522098
rect 67408 521778 67450 522014
rect 67686 521778 67728 522014
rect 67408 521746 67728 521778
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 62288 482614 62608 482646
rect 62288 482378 62330 482614
rect 62566 482378 62608 482614
rect 62288 482294 62608 482378
rect 62288 482058 62330 482294
rect 62566 482058 62608 482294
rect 62288 482026 62608 482058
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 57168 442894 57488 442926
rect 57168 442658 57210 442894
rect 57446 442658 57488 442894
rect 57168 442574 57488 442658
rect 57168 442338 57210 442574
rect 57446 442338 57488 442574
rect 57168 442306 57488 442338
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 60114 421774 60734 457218
rect 63834 461494 64454 496938
rect 73794 507454 74414 542898
rect 77648 543454 77968 543486
rect 77648 543218 77690 543454
rect 77926 543218 77968 543454
rect 77648 543134 77968 543218
rect 77648 542898 77690 543134
rect 77926 542898 77968 543134
rect 77648 542866 77968 542898
rect 81234 514894 81854 550338
rect 84954 554614 85574 590058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 630334 89294 665778
rect 88674 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 89294 630334
rect 88674 630014 89294 630098
rect 88674 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 89294 630014
rect 88674 594334 89294 629778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 602500 93014 633498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 88674 594098 88706 594334
rect 88942 594098 89026 594334
rect 89262 594098 89294 594334
rect 88674 594014 89294 594098
rect 88674 593778 88706 594014
rect 88942 593778 89026 594014
rect 89262 593778 89294 594014
rect 87888 586894 88208 586926
rect 87888 586658 87930 586894
rect 88166 586658 88208 586894
rect 87888 586574 88208 586658
rect 87888 586338 87930 586574
rect 88166 586338 88208 586574
rect 87888 586306 88208 586338
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 82768 547174 83088 547206
rect 82768 546938 82810 547174
rect 83046 546938 83088 547174
rect 82768 546854 83088 546938
rect 82768 546618 82810 546854
rect 83046 546618 83088 546854
rect 82768 546586 83088 546618
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 72528 490054 72848 490086
rect 72528 489818 72570 490054
rect 72806 489818 72848 490054
rect 72528 489734 72848 489818
rect 72528 489498 72570 489734
rect 72806 489498 72848 489734
rect 72528 489466 72848 489498
rect 67408 486334 67728 486366
rect 67408 486098 67450 486334
rect 67686 486098 67728 486334
rect 67408 486014 67728 486098
rect 67408 485778 67450 486014
rect 67686 485778 67728 486014
rect 67408 485746 67728 485778
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 62288 446614 62608 446646
rect 62288 446378 62330 446614
rect 62566 446378 62608 446614
rect 62288 446294 62608 446378
rect 62288 446058 62330 446294
rect 62566 446058 62608 446294
rect 62288 446026 62608 446058
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 57168 406894 57488 406926
rect 57168 406658 57210 406894
rect 57446 406658 57488 406894
rect 57168 406574 57488 406658
rect 57168 406338 57210 406574
rect 57446 406338 57488 406574
rect 57168 406306 57488 406338
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 60114 385774 60734 421218
rect 63834 425494 64454 460938
rect 73794 471454 74414 506898
rect 77648 507454 77968 507486
rect 77648 507218 77690 507454
rect 77926 507218 77968 507454
rect 77648 507134 77968 507218
rect 77648 506898 77690 507134
rect 77926 506898 77968 507134
rect 77648 506866 77968 506898
rect 81234 478894 81854 514338
rect 84954 518614 85574 554058
rect 88674 558334 89294 593778
rect 96114 601774 96734 637218
rect 96114 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 96734 601774
rect 96114 601454 96734 601538
rect 96114 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 96734 601454
rect 93008 590614 93328 590646
rect 93008 590378 93050 590614
rect 93286 590378 93328 590614
rect 93008 590294 93328 590378
rect 93008 590058 93050 590294
rect 93286 590058 93328 590294
rect 93008 590026 93328 590058
rect 88674 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 89294 558334
rect 88674 558014 89294 558098
rect 88674 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 89294 558014
rect 87888 550894 88208 550926
rect 87888 550658 87930 550894
rect 88166 550658 88208 550894
rect 87888 550574 88208 550658
rect 87888 550338 87930 550574
rect 88166 550338 88208 550574
rect 87888 550306 88208 550338
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 82768 511174 83088 511206
rect 82768 510938 82810 511174
rect 83046 510938 83088 511174
rect 82768 510854 83088 510938
rect 82768 510618 82810 510854
rect 83046 510618 83088 510854
rect 82768 510586 83088 510618
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 72528 454054 72848 454086
rect 72528 453818 72570 454054
rect 72806 453818 72848 454054
rect 72528 453734 72848 453818
rect 72528 453498 72570 453734
rect 72806 453498 72848 453734
rect 72528 453466 72848 453498
rect 67408 450334 67728 450366
rect 67408 450098 67450 450334
rect 67686 450098 67728 450334
rect 67408 450014 67728 450098
rect 67408 449778 67450 450014
rect 67686 449778 67728 450014
rect 67408 449746 67728 449778
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 62288 410614 62608 410646
rect 62288 410378 62330 410614
rect 62566 410378 62608 410614
rect 62288 410294 62608 410378
rect 62288 410058 62330 410294
rect 62566 410058 62608 410294
rect 62288 410026 62608 410058
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 57168 370894 57488 370926
rect 57168 370658 57210 370894
rect 57446 370658 57488 370894
rect 57168 370574 57488 370658
rect 57168 370338 57210 370574
rect 57446 370338 57488 370574
rect 57168 370306 57488 370338
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 60114 349774 60734 385218
rect 63834 389494 64454 424938
rect 73794 435454 74414 470898
rect 77648 471454 77968 471486
rect 77648 471218 77690 471454
rect 77926 471218 77968 471454
rect 77648 471134 77968 471218
rect 77648 470898 77690 471134
rect 77926 470898 77968 471134
rect 77648 470866 77968 470898
rect 81234 442894 81854 478338
rect 84954 482614 85574 518058
rect 88674 522334 89294 557778
rect 96114 565774 96734 601218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 605494 100454 640938
rect 99834 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 100454 605494
rect 99834 605174 100454 605258
rect 99834 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 100454 605174
rect 98128 594334 98448 594366
rect 98128 594098 98170 594334
rect 98406 594098 98448 594334
rect 98128 594014 98448 594098
rect 98128 593778 98170 594014
rect 98406 593778 98448 594014
rect 98128 593746 98448 593778
rect 96114 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 96734 565774
rect 96114 565454 96734 565538
rect 96114 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 96734 565454
rect 93008 554614 93328 554646
rect 93008 554378 93050 554614
rect 93286 554378 93328 554614
rect 93008 554294 93328 554378
rect 93008 554058 93050 554294
rect 93286 554058 93328 554294
rect 93008 554026 93328 554058
rect 88674 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 89294 522334
rect 88674 522014 89294 522098
rect 88674 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 89294 522014
rect 87888 514894 88208 514926
rect 87888 514658 87930 514894
rect 88166 514658 88208 514894
rect 87888 514574 88208 514658
rect 87888 514338 87930 514574
rect 88166 514338 88208 514574
rect 87888 514306 88208 514338
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 82768 475174 83088 475206
rect 82768 474938 82810 475174
rect 83046 474938 83088 475174
rect 82768 474854 83088 474938
rect 82768 474618 82810 474854
rect 83046 474618 83088 474854
rect 82768 474586 83088 474618
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 72528 418054 72848 418086
rect 72528 417818 72570 418054
rect 72806 417818 72848 418054
rect 72528 417734 72848 417818
rect 72528 417498 72570 417734
rect 72806 417498 72848 417734
rect 72528 417466 72848 417498
rect 67408 414334 67728 414366
rect 67408 414098 67450 414334
rect 67686 414098 67728 414334
rect 67408 414014 67728 414098
rect 67408 413778 67450 414014
rect 67686 413778 67728 414014
rect 67408 413746 67728 413778
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 62288 374614 62608 374646
rect 62288 374378 62330 374614
rect 62566 374378 62608 374614
rect 62288 374294 62608 374378
rect 62288 374058 62330 374294
rect 62566 374058 62608 374294
rect 62288 374026 62608 374058
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 57168 334894 57488 334926
rect 57168 334658 57210 334894
rect 57446 334658 57488 334894
rect 57168 334574 57488 334658
rect 57168 334338 57210 334574
rect 57446 334338 57488 334574
rect 57168 334306 57488 334338
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 60114 313774 60734 349218
rect 63834 353494 64454 388938
rect 73794 399454 74414 434898
rect 77648 435454 77968 435486
rect 77648 435218 77690 435454
rect 77926 435218 77968 435454
rect 77648 435134 77968 435218
rect 77648 434898 77690 435134
rect 77926 434898 77968 435134
rect 77648 434866 77968 434898
rect 81234 406894 81854 442338
rect 84954 446614 85574 482058
rect 88674 486334 89294 521778
rect 96114 529774 96734 565218
rect 99834 569494 100454 604938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 103248 598054 103568 598086
rect 103248 597818 103290 598054
rect 103526 597818 103568 598054
rect 103248 597734 103568 597818
rect 103248 597498 103290 597734
rect 103526 597498 103568 597734
rect 103248 597466 103568 597498
rect 108368 579454 108688 579486
rect 108368 579218 108410 579454
rect 108646 579218 108688 579454
rect 108368 579134 108688 579218
rect 108368 578898 108410 579134
rect 108646 578898 108688 579134
rect 108368 578866 108688 578898
rect 109794 579454 110414 614898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 602500 114134 618618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 630334 125294 665778
rect 124674 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 125294 630334
rect 124674 630014 125294 630098
rect 124674 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 125294 630014
rect 124674 594334 125294 629778
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 602500 129014 633498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 601774 132734 637218
rect 132114 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 132734 601774
rect 132114 601454 132734 601538
rect 132114 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 132734 601454
rect 124674 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 125294 594334
rect 124674 594014 125294 594098
rect 124674 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 125294 594014
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 113488 583174 113808 583206
rect 113488 582938 113530 583174
rect 113766 582938 113808 583174
rect 113488 582854 113808 582938
rect 113488 582618 113530 582854
rect 113766 582618 113808 582854
rect 113488 582586 113808 582618
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 99834 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 100454 569494
rect 99834 569174 100454 569258
rect 99834 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 100454 569174
rect 98128 558334 98448 558366
rect 98128 558098 98170 558334
rect 98406 558098 98448 558334
rect 98128 558014 98448 558098
rect 98128 557778 98170 558014
rect 98406 557778 98448 558014
rect 98128 557746 98448 557778
rect 96114 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 96734 529774
rect 96114 529454 96734 529538
rect 96114 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 96734 529454
rect 93008 518614 93328 518646
rect 93008 518378 93050 518614
rect 93286 518378 93328 518614
rect 93008 518294 93328 518378
rect 93008 518058 93050 518294
rect 93286 518058 93328 518294
rect 93008 518026 93328 518058
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 87888 478894 88208 478926
rect 87888 478658 87930 478894
rect 88166 478658 88208 478894
rect 87888 478574 88208 478658
rect 87888 478338 87930 478574
rect 88166 478338 88208 478574
rect 87888 478306 88208 478338
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 82768 439174 83088 439206
rect 82768 438938 82810 439174
rect 83046 438938 83088 439174
rect 82768 438854 83088 438938
rect 82768 438618 82810 438854
rect 83046 438618 83088 438854
rect 82768 438586 83088 438618
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 72528 382054 72848 382086
rect 72528 381818 72570 382054
rect 72806 381818 72848 382054
rect 72528 381734 72848 381818
rect 72528 381498 72570 381734
rect 72806 381498 72848 381734
rect 72528 381466 72848 381498
rect 67408 378334 67728 378366
rect 67408 378098 67450 378334
rect 67686 378098 67728 378334
rect 67408 378014 67728 378098
rect 67408 377778 67450 378014
rect 67686 377778 67728 378014
rect 67408 377746 67728 377778
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 62288 338614 62608 338646
rect 62288 338378 62330 338614
rect 62566 338378 62608 338614
rect 62288 338294 62608 338378
rect 62288 338058 62330 338294
rect 62566 338058 62608 338294
rect 62288 338026 62608 338058
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 57168 298894 57488 298926
rect 57168 298658 57210 298894
rect 57446 298658 57488 298894
rect 57168 298574 57488 298658
rect 57168 298338 57210 298574
rect 57446 298338 57488 298574
rect 57168 298306 57488 298338
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 60114 277774 60734 313218
rect 63834 317494 64454 352938
rect 73794 363454 74414 398898
rect 77648 399454 77968 399486
rect 77648 399218 77690 399454
rect 77926 399218 77968 399454
rect 77648 399134 77968 399218
rect 77648 398898 77690 399134
rect 77926 398898 77968 399134
rect 77648 398866 77968 398898
rect 81234 370894 81854 406338
rect 84954 410614 85574 446058
rect 88674 450334 89294 485778
rect 96114 493774 96734 529218
rect 99834 533494 100454 568938
rect 103248 562054 103568 562086
rect 103248 561818 103290 562054
rect 103526 561818 103568 562054
rect 103248 561734 103568 561818
rect 103248 561498 103290 561734
rect 103526 561498 103568 561734
rect 103248 561466 103568 561498
rect 108368 543454 108688 543486
rect 108368 543218 108410 543454
rect 108646 543218 108688 543454
rect 108368 543134 108688 543218
rect 108368 542898 108410 543134
rect 108646 542898 108688 543134
rect 108368 542866 108688 542898
rect 109794 543454 110414 578898
rect 117234 550894 117854 586338
rect 118608 586894 118928 586926
rect 118608 586658 118650 586894
rect 118886 586658 118928 586894
rect 118608 586574 118928 586658
rect 118608 586338 118650 586574
rect 118886 586338 118928 586574
rect 118608 586306 118928 586338
rect 120954 554614 121574 590058
rect 123728 590614 124048 590646
rect 123728 590378 123770 590614
rect 124006 590378 124048 590614
rect 123728 590294 124048 590378
rect 123728 590058 123770 590294
rect 124006 590058 124048 590294
rect 123728 590026 124048 590058
rect 124674 558334 125294 593778
rect 128848 594334 129168 594366
rect 128848 594098 128890 594334
rect 129126 594098 129168 594334
rect 128848 594014 129168 594098
rect 128848 593778 128890 594014
rect 129126 593778 129168 594014
rect 128848 593746 129168 593778
rect 132114 565774 132734 601218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 135834 605494 136454 640938
rect 135834 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 136454 605494
rect 135834 605174 136454 605258
rect 135834 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 136454 605174
rect 133968 598054 134288 598086
rect 133968 597818 134010 598054
rect 134246 597818 134288 598054
rect 133968 597734 134288 597818
rect 133968 597498 134010 597734
rect 134246 597498 134288 597734
rect 133968 597466 134288 597498
rect 132114 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 132734 565774
rect 132114 565454 132734 565538
rect 132114 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 132734 565454
rect 124674 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 125294 558334
rect 124674 558014 125294 558098
rect 124674 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 125294 558014
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 113488 547174 113808 547206
rect 113488 546938 113530 547174
rect 113766 546938 113808 547174
rect 113488 546854 113808 546938
rect 113488 546618 113530 546854
rect 113766 546618 113808 546854
rect 113488 546586 113808 546618
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 99834 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 100454 533494
rect 99834 533174 100454 533258
rect 99834 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 100454 533174
rect 98128 522334 98448 522366
rect 98128 522098 98170 522334
rect 98406 522098 98448 522334
rect 98128 522014 98448 522098
rect 98128 521778 98170 522014
rect 98406 521778 98448 522014
rect 98128 521746 98448 521778
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 93008 482614 93328 482646
rect 93008 482378 93050 482614
rect 93286 482378 93328 482614
rect 93008 482294 93328 482378
rect 93008 482058 93050 482294
rect 93286 482058 93328 482294
rect 93008 482026 93328 482058
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 87888 442894 88208 442926
rect 87888 442658 87930 442894
rect 88166 442658 88208 442894
rect 87888 442574 88208 442658
rect 87888 442338 87930 442574
rect 88166 442338 88208 442574
rect 87888 442306 88208 442338
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 82768 403174 83088 403206
rect 82768 402938 82810 403174
rect 83046 402938 83088 403174
rect 82768 402854 83088 402938
rect 82768 402618 82810 402854
rect 83046 402618 83088 402854
rect 82768 402586 83088 402618
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 72528 346054 72848 346086
rect 72528 345818 72570 346054
rect 72806 345818 72848 346054
rect 72528 345734 72848 345818
rect 72528 345498 72570 345734
rect 72806 345498 72848 345734
rect 72528 345466 72848 345498
rect 67408 342334 67728 342366
rect 67408 342098 67450 342334
rect 67686 342098 67728 342334
rect 67408 342014 67728 342098
rect 67408 341778 67450 342014
rect 67686 341778 67728 342014
rect 67408 341746 67728 341778
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 62288 302614 62608 302646
rect 62288 302378 62330 302614
rect 62566 302378 62608 302614
rect 62288 302294 62608 302378
rect 62288 302058 62330 302294
rect 62566 302058 62608 302294
rect 62288 302026 62608 302058
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 57168 262894 57488 262926
rect 57168 262658 57210 262894
rect 57446 262658 57488 262894
rect 57168 262574 57488 262658
rect 57168 262338 57210 262574
rect 57446 262338 57488 262574
rect 57168 262306 57488 262338
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 60114 241774 60734 277218
rect 63834 281494 64454 316938
rect 73794 327454 74414 362898
rect 77648 363454 77968 363486
rect 77648 363218 77690 363454
rect 77926 363218 77968 363454
rect 77648 363134 77968 363218
rect 77648 362898 77690 363134
rect 77926 362898 77968 363134
rect 77648 362866 77968 362898
rect 81234 334894 81854 370338
rect 84954 374614 85574 410058
rect 88674 414334 89294 449778
rect 96114 457774 96734 493218
rect 99834 497494 100454 532938
rect 103248 526054 103568 526086
rect 103248 525818 103290 526054
rect 103526 525818 103568 526054
rect 103248 525734 103568 525818
rect 103248 525498 103290 525734
rect 103526 525498 103568 525734
rect 103248 525466 103568 525498
rect 108368 507454 108688 507486
rect 108368 507218 108410 507454
rect 108646 507218 108688 507454
rect 108368 507134 108688 507218
rect 108368 506898 108410 507134
rect 108646 506898 108688 507134
rect 108368 506866 108688 506898
rect 109794 507454 110414 542898
rect 117234 514894 117854 550338
rect 118608 550894 118928 550926
rect 118608 550658 118650 550894
rect 118886 550658 118928 550894
rect 118608 550574 118928 550658
rect 118608 550338 118650 550574
rect 118886 550338 118928 550574
rect 118608 550306 118928 550338
rect 120954 518614 121574 554058
rect 123728 554614 124048 554646
rect 123728 554378 123770 554614
rect 124006 554378 124048 554614
rect 123728 554294 124048 554378
rect 123728 554058 123770 554294
rect 124006 554058 124048 554294
rect 123728 554026 124048 554058
rect 124674 522334 125294 557778
rect 128848 558334 129168 558366
rect 128848 558098 128890 558334
rect 129126 558098 129168 558334
rect 128848 558014 129168 558098
rect 128848 557778 128890 558014
rect 129126 557778 129168 558014
rect 128848 557746 129168 557778
rect 132114 529774 132734 565218
rect 135834 569494 136454 604938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 144208 583174 144528 583206
rect 144208 582938 144250 583174
rect 144486 582938 144528 583174
rect 144208 582854 144528 582938
rect 144208 582618 144250 582854
rect 144486 582618 144528 582854
rect 144208 582586 144528 582618
rect 139088 579454 139408 579486
rect 139088 579218 139130 579454
rect 139366 579218 139408 579454
rect 139088 579134 139408 579218
rect 139088 578898 139130 579134
rect 139366 578898 139408 579134
rect 139088 578866 139408 578898
rect 145794 579454 146414 614898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 602500 150134 618618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 149328 586894 149648 586926
rect 149328 586658 149370 586894
rect 149606 586658 149648 586894
rect 149328 586574 149648 586658
rect 149328 586338 149370 586574
rect 149606 586338 149648 586574
rect 149328 586306 149648 586338
rect 153234 586894 153854 622338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 154448 590614 154768 590646
rect 154448 590378 154490 590614
rect 154726 590378 154768 590614
rect 154448 590294 154768 590378
rect 154448 590058 154490 590294
rect 154726 590058 154768 590294
rect 154448 590026 154768 590058
rect 156954 590614 157574 626058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 159568 594334 159888 594366
rect 159568 594098 159610 594334
rect 159846 594098 159888 594334
rect 159568 594014 159888 594098
rect 159568 593778 159610 594014
rect 159846 593778 159888 594014
rect 159568 593746 159888 593778
rect 160674 594334 161294 629778
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 602500 165014 633498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 164688 598054 165008 598086
rect 164688 597818 164730 598054
rect 164966 597818 165008 598054
rect 164688 597734 165008 597818
rect 164688 597498 164730 597734
rect 164966 597498 165008 597734
rect 164688 597466 165008 597498
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 135834 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 136454 569494
rect 135834 569174 136454 569258
rect 135834 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 136454 569174
rect 133968 562054 134288 562086
rect 133968 561818 134010 562054
rect 134246 561818 134288 562054
rect 133968 561734 134288 561818
rect 133968 561498 134010 561734
rect 134246 561498 134288 561734
rect 133968 561466 134288 561498
rect 132114 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 132734 529774
rect 132114 529454 132734 529538
rect 132114 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 132734 529454
rect 124674 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 125294 522334
rect 124674 522014 125294 522098
rect 124674 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 125294 522014
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 113488 511174 113808 511206
rect 113488 510938 113530 511174
rect 113766 510938 113808 511174
rect 113488 510854 113808 510938
rect 113488 510618 113530 510854
rect 113766 510618 113808 510854
rect 113488 510586 113808 510618
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 98128 486334 98448 486366
rect 98128 486098 98170 486334
rect 98406 486098 98448 486334
rect 98128 486014 98448 486098
rect 98128 485778 98170 486014
rect 98406 485778 98448 486014
rect 98128 485746 98448 485778
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 93008 446614 93328 446646
rect 93008 446378 93050 446614
rect 93286 446378 93328 446614
rect 93008 446294 93328 446378
rect 93008 446058 93050 446294
rect 93286 446058 93328 446294
rect 93008 446026 93328 446058
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 87888 406894 88208 406926
rect 87888 406658 87930 406894
rect 88166 406658 88208 406894
rect 87888 406574 88208 406658
rect 87888 406338 87930 406574
rect 88166 406338 88208 406574
rect 87888 406306 88208 406338
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 82768 367174 83088 367206
rect 82768 366938 82810 367174
rect 83046 366938 83088 367174
rect 82768 366854 83088 366938
rect 82768 366618 82810 366854
rect 83046 366618 83088 366854
rect 82768 366586 83088 366618
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 72528 310054 72848 310086
rect 72528 309818 72570 310054
rect 72806 309818 72848 310054
rect 72528 309734 72848 309818
rect 72528 309498 72570 309734
rect 72806 309498 72848 309734
rect 72528 309466 72848 309498
rect 67408 306334 67728 306366
rect 67408 306098 67450 306334
rect 67686 306098 67728 306334
rect 67408 306014 67728 306098
rect 67408 305778 67450 306014
rect 67686 305778 67728 306014
rect 67408 305746 67728 305778
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 62288 266614 62608 266646
rect 62288 266378 62330 266614
rect 62566 266378 62608 266614
rect 62288 266294 62608 266378
rect 62288 266058 62330 266294
rect 62566 266058 62608 266294
rect 62288 266026 62608 266058
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 57168 226894 57488 226926
rect 57168 226658 57210 226894
rect 57446 226658 57488 226894
rect 57168 226574 57488 226658
rect 57168 226338 57210 226574
rect 57446 226338 57488 226574
rect 57168 226306 57488 226338
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 60114 205774 60734 241218
rect 63834 245494 64454 280938
rect 73794 291454 74414 326898
rect 77648 327454 77968 327486
rect 77648 327218 77690 327454
rect 77926 327218 77968 327454
rect 77648 327134 77968 327218
rect 77648 326898 77690 327134
rect 77926 326898 77968 327134
rect 77648 326866 77968 326898
rect 81234 298894 81854 334338
rect 84954 338614 85574 374058
rect 88674 378334 89294 413778
rect 96114 421774 96734 457218
rect 99834 461494 100454 496938
rect 103248 490054 103568 490086
rect 103248 489818 103290 490054
rect 103526 489818 103568 490054
rect 103248 489734 103568 489818
rect 103248 489498 103290 489734
rect 103526 489498 103568 489734
rect 103248 489466 103568 489498
rect 108368 471454 108688 471486
rect 108368 471218 108410 471454
rect 108646 471218 108688 471454
rect 108368 471134 108688 471218
rect 108368 470898 108410 471134
rect 108646 470898 108688 471134
rect 108368 470866 108688 470898
rect 109794 471454 110414 506898
rect 117234 478894 117854 514338
rect 118608 514894 118928 514926
rect 118608 514658 118650 514894
rect 118886 514658 118928 514894
rect 118608 514574 118928 514658
rect 118608 514338 118650 514574
rect 118886 514338 118928 514574
rect 118608 514306 118928 514338
rect 120954 482614 121574 518058
rect 123728 518614 124048 518646
rect 123728 518378 123770 518614
rect 124006 518378 124048 518614
rect 123728 518294 124048 518378
rect 123728 518058 123770 518294
rect 124006 518058 124048 518294
rect 123728 518026 124048 518058
rect 124674 486334 125294 521778
rect 128848 522334 129168 522366
rect 128848 522098 128890 522334
rect 129126 522098 129168 522334
rect 128848 522014 129168 522098
rect 128848 521778 128890 522014
rect 129126 521778 129168 522014
rect 128848 521746 129168 521778
rect 132114 493774 132734 529218
rect 135834 533494 136454 568938
rect 144208 547174 144528 547206
rect 144208 546938 144250 547174
rect 144486 546938 144528 547174
rect 144208 546854 144528 546938
rect 144208 546618 144250 546854
rect 144486 546618 144528 546854
rect 144208 546586 144528 546618
rect 139088 543454 139408 543486
rect 139088 543218 139130 543454
rect 139366 543218 139408 543454
rect 139088 543134 139408 543218
rect 139088 542898 139130 543134
rect 139366 542898 139408 543134
rect 139088 542866 139408 542898
rect 145794 543454 146414 578898
rect 149328 550894 149648 550926
rect 149328 550658 149370 550894
rect 149606 550658 149648 550894
rect 149328 550574 149648 550658
rect 149328 550338 149370 550574
rect 149606 550338 149648 550574
rect 149328 550306 149648 550338
rect 153234 550894 153854 586338
rect 154448 554614 154768 554646
rect 154448 554378 154490 554614
rect 154726 554378 154768 554614
rect 154448 554294 154768 554378
rect 154448 554058 154490 554294
rect 154726 554058 154768 554294
rect 154448 554026 154768 554058
rect 156954 554614 157574 590058
rect 159568 558334 159888 558366
rect 159568 558098 159610 558334
rect 159846 558098 159888 558334
rect 159568 558014 159888 558098
rect 159568 557778 159610 558014
rect 159846 557778 159888 558014
rect 159568 557746 159888 557778
rect 160674 558334 161294 593778
rect 168114 565774 168734 601218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 169808 579454 170128 579486
rect 169808 579218 169850 579454
rect 170086 579218 170128 579454
rect 169808 579134 170128 579218
rect 169808 578898 169850 579134
rect 170086 578898 170128 579134
rect 169808 578866 170128 578898
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 164688 562054 165008 562086
rect 164688 561818 164730 562054
rect 164966 561818 165008 562054
rect 164688 561734 165008 561818
rect 164688 561498 164730 561734
rect 164966 561498 165008 561734
rect 164688 561466 165008 561498
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 135834 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 136454 533494
rect 135834 533174 136454 533258
rect 135834 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 136454 533174
rect 133968 526054 134288 526086
rect 133968 525818 134010 526054
rect 134246 525818 134288 526054
rect 133968 525734 134288 525818
rect 133968 525498 134010 525734
rect 134246 525498 134288 525734
rect 133968 525466 134288 525498
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 113488 475174 113808 475206
rect 113488 474938 113530 475174
rect 113766 474938 113808 475174
rect 113488 474854 113808 474938
rect 113488 474618 113530 474854
rect 113766 474618 113808 474854
rect 113488 474586 113808 474618
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 98128 450334 98448 450366
rect 98128 450098 98170 450334
rect 98406 450098 98448 450334
rect 98128 450014 98448 450098
rect 98128 449778 98170 450014
rect 98406 449778 98448 450014
rect 98128 449746 98448 449778
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 93008 410614 93328 410646
rect 93008 410378 93050 410614
rect 93286 410378 93328 410614
rect 93008 410294 93328 410378
rect 93008 410058 93050 410294
rect 93286 410058 93328 410294
rect 93008 410026 93328 410058
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 87888 370894 88208 370926
rect 87888 370658 87930 370894
rect 88166 370658 88208 370894
rect 87888 370574 88208 370658
rect 87888 370338 87930 370574
rect 88166 370338 88208 370574
rect 87888 370306 88208 370338
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 82768 331174 83088 331206
rect 82768 330938 82810 331174
rect 83046 330938 83088 331174
rect 82768 330854 83088 330938
rect 82768 330618 82810 330854
rect 83046 330618 83088 330854
rect 82768 330586 83088 330618
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 72528 274054 72848 274086
rect 72528 273818 72570 274054
rect 72806 273818 72848 274054
rect 72528 273734 72848 273818
rect 72528 273498 72570 273734
rect 72806 273498 72848 273734
rect 72528 273466 72848 273498
rect 67408 270334 67728 270366
rect 67408 270098 67450 270334
rect 67686 270098 67728 270334
rect 67408 270014 67728 270098
rect 67408 269778 67450 270014
rect 67686 269778 67728 270014
rect 67408 269746 67728 269778
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 62288 230614 62608 230646
rect 62288 230378 62330 230614
rect 62566 230378 62608 230614
rect 62288 230294 62608 230378
rect 62288 230058 62330 230294
rect 62566 230058 62608 230294
rect 62288 230026 62608 230058
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 57168 190894 57488 190926
rect 57168 190658 57210 190894
rect 57446 190658 57488 190894
rect 57168 190574 57488 190658
rect 57168 190338 57210 190574
rect 57446 190338 57488 190574
rect 57168 190306 57488 190338
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 130054 57014 165498
rect 60114 169774 60734 205218
rect 63834 209494 64454 244938
rect 73794 255454 74414 290898
rect 77648 291454 77968 291486
rect 77648 291218 77690 291454
rect 77926 291218 77968 291454
rect 77648 291134 77968 291218
rect 77648 290898 77690 291134
rect 77926 290898 77968 291134
rect 77648 290866 77968 290898
rect 81234 262894 81854 298338
rect 84954 302614 85574 338058
rect 88674 342334 89294 377778
rect 96114 385774 96734 421218
rect 99834 425494 100454 460938
rect 103248 454054 103568 454086
rect 103248 453818 103290 454054
rect 103526 453818 103568 454054
rect 103248 453734 103568 453818
rect 103248 453498 103290 453734
rect 103526 453498 103568 453734
rect 103248 453466 103568 453498
rect 108368 435454 108688 435486
rect 108368 435218 108410 435454
rect 108646 435218 108688 435454
rect 108368 435134 108688 435218
rect 108368 434898 108410 435134
rect 108646 434898 108688 435134
rect 108368 434866 108688 434898
rect 109794 435454 110414 470898
rect 117234 442894 117854 478338
rect 118608 478894 118928 478926
rect 118608 478658 118650 478894
rect 118886 478658 118928 478894
rect 118608 478574 118928 478658
rect 118608 478338 118650 478574
rect 118886 478338 118928 478574
rect 118608 478306 118928 478338
rect 120954 446614 121574 482058
rect 123728 482614 124048 482646
rect 123728 482378 123770 482614
rect 124006 482378 124048 482614
rect 123728 482294 124048 482378
rect 123728 482058 123770 482294
rect 124006 482058 124048 482294
rect 123728 482026 124048 482058
rect 124674 450334 125294 485778
rect 128848 486334 129168 486366
rect 128848 486098 128890 486334
rect 129126 486098 129168 486334
rect 128848 486014 129168 486098
rect 128848 485778 128890 486014
rect 129126 485778 129168 486014
rect 128848 485746 129168 485778
rect 132114 457774 132734 493218
rect 135834 497494 136454 532938
rect 144208 511174 144528 511206
rect 144208 510938 144250 511174
rect 144486 510938 144528 511174
rect 144208 510854 144528 510938
rect 144208 510618 144250 510854
rect 144486 510618 144528 510854
rect 144208 510586 144528 510618
rect 139088 507454 139408 507486
rect 139088 507218 139130 507454
rect 139366 507218 139408 507454
rect 139088 507134 139408 507218
rect 139088 506898 139130 507134
rect 139366 506898 139408 507134
rect 139088 506866 139408 506898
rect 145794 507454 146414 542898
rect 149328 514894 149648 514926
rect 149328 514658 149370 514894
rect 149606 514658 149648 514894
rect 149328 514574 149648 514658
rect 149328 514338 149370 514574
rect 149606 514338 149648 514574
rect 149328 514306 149648 514338
rect 153234 514894 153854 550338
rect 154448 518614 154768 518646
rect 154448 518378 154490 518614
rect 154726 518378 154768 518614
rect 154448 518294 154768 518378
rect 154448 518058 154490 518294
rect 154726 518058 154768 518294
rect 154448 518026 154768 518058
rect 156954 518614 157574 554058
rect 159568 522334 159888 522366
rect 159568 522098 159610 522334
rect 159846 522098 159888 522334
rect 159568 522014 159888 522098
rect 159568 521778 159610 522014
rect 159846 521778 159888 522014
rect 159568 521746 159888 521778
rect 160674 522334 161294 557778
rect 168114 529774 168734 565218
rect 171834 569494 172454 604938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 180048 586894 180368 586926
rect 180048 586658 180090 586894
rect 180326 586658 180368 586894
rect 180048 586574 180368 586658
rect 180048 586338 180090 586574
rect 180326 586338 180368 586574
rect 180048 586306 180368 586338
rect 174928 583174 175248 583206
rect 174928 582938 174970 583174
rect 175206 582938 175248 583174
rect 174928 582854 175248 582938
rect 174928 582618 174970 582854
rect 175206 582618 175248 582854
rect 174928 582586 175248 582618
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 169808 543454 170128 543486
rect 169808 543218 169850 543454
rect 170086 543218 170128 543454
rect 169808 543134 170128 543218
rect 169808 542898 169850 543134
rect 170086 542898 170128 543134
rect 169808 542866 170128 542898
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 164688 526054 165008 526086
rect 164688 525818 164730 526054
rect 164966 525818 165008 526054
rect 164688 525734 165008 525818
rect 164688 525498 164730 525734
rect 164966 525498 165008 525734
rect 164688 525466 165008 525498
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 133968 490054 134288 490086
rect 133968 489818 134010 490054
rect 134246 489818 134288 490054
rect 133968 489734 134288 489818
rect 133968 489498 134010 489734
rect 134246 489498 134288 489734
rect 133968 489466 134288 489498
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 113488 439174 113808 439206
rect 113488 438938 113530 439174
rect 113766 438938 113808 439174
rect 113488 438854 113808 438938
rect 113488 438618 113530 438854
rect 113766 438618 113808 438854
rect 113488 438586 113808 438618
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 98128 414334 98448 414366
rect 98128 414098 98170 414334
rect 98406 414098 98448 414334
rect 98128 414014 98448 414098
rect 98128 413778 98170 414014
rect 98406 413778 98448 414014
rect 98128 413746 98448 413778
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 93008 374614 93328 374646
rect 93008 374378 93050 374614
rect 93286 374378 93328 374614
rect 93008 374294 93328 374378
rect 93008 374058 93050 374294
rect 93286 374058 93328 374294
rect 93008 374026 93328 374058
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 87888 334894 88208 334926
rect 87888 334658 87930 334894
rect 88166 334658 88208 334894
rect 87888 334574 88208 334658
rect 87888 334338 87930 334574
rect 88166 334338 88208 334574
rect 87888 334306 88208 334338
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 82768 295174 83088 295206
rect 82768 294938 82810 295174
rect 83046 294938 83088 295174
rect 82768 294854 83088 294938
rect 82768 294618 82810 294854
rect 83046 294618 83088 294854
rect 82768 294586 83088 294618
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 72528 238054 72848 238086
rect 72528 237818 72570 238054
rect 72806 237818 72848 238054
rect 72528 237734 72848 237818
rect 72528 237498 72570 237734
rect 72806 237498 72848 237734
rect 72528 237466 72848 237498
rect 67408 234334 67728 234366
rect 67408 234098 67450 234334
rect 67686 234098 67728 234334
rect 67408 234014 67728 234098
rect 67408 233778 67450 234014
rect 67686 233778 67728 234014
rect 67408 233746 67728 233778
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 62288 194614 62608 194646
rect 62288 194378 62330 194614
rect 62566 194378 62608 194614
rect 62288 194294 62608 194378
rect 62288 194058 62330 194294
rect 62566 194058 62608 194294
rect 62288 194026 62608 194058
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 57168 154894 57488 154926
rect 57168 154658 57210 154894
rect 57446 154658 57488 154894
rect 57168 154574 57488 154658
rect 57168 154338 57210 154574
rect 57446 154338 57488 154574
rect 57168 154306 57488 154338
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 56394 94054 57014 129498
rect 60114 133774 60734 169218
rect 63834 173494 64454 208938
rect 73794 219454 74414 254898
rect 77648 255454 77968 255486
rect 77648 255218 77690 255454
rect 77926 255218 77968 255454
rect 77648 255134 77968 255218
rect 77648 254898 77690 255134
rect 77926 254898 77968 255134
rect 77648 254866 77968 254898
rect 81234 226894 81854 262338
rect 84954 266614 85574 302058
rect 88674 306334 89294 341778
rect 96114 349774 96734 385218
rect 99834 389494 100454 424938
rect 103248 418054 103568 418086
rect 103248 417818 103290 418054
rect 103526 417818 103568 418054
rect 103248 417734 103568 417818
rect 103248 417498 103290 417734
rect 103526 417498 103568 417734
rect 103248 417466 103568 417498
rect 108368 399454 108688 399486
rect 108368 399218 108410 399454
rect 108646 399218 108688 399454
rect 108368 399134 108688 399218
rect 108368 398898 108410 399134
rect 108646 398898 108688 399134
rect 108368 398866 108688 398898
rect 109794 399454 110414 434898
rect 117234 406894 117854 442338
rect 118608 442894 118928 442926
rect 118608 442658 118650 442894
rect 118886 442658 118928 442894
rect 118608 442574 118928 442658
rect 118608 442338 118650 442574
rect 118886 442338 118928 442574
rect 118608 442306 118928 442338
rect 120954 410614 121574 446058
rect 123728 446614 124048 446646
rect 123728 446378 123770 446614
rect 124006 446378 124048 446614
rect 123728 446294 124048 446378
rect 123728 446058 123770 446294
rect 124006 446058 124048 446294
rect 123728 446026 124048 446058
rect 124674 414334 125294 449778
rect 128848 450334 129168 450366
rect 128848 450098 128890 450334
rect 129126 450098 129168 450334
rect 128848 450014 129168 450098
rect 128848 449778 128890 450014
rect 129126 449778 129168 450014
rect 128848 449746 129168 449778
rect 132114 421774 132734 457218
rect 135834 461494 136454 496938
rect 144208 475174 144528 475206
rect 144208 474938 144250 475174
rect 144486 474938 144528 475174
rect 144208 474854 144528 474938
rect 144208 474618 144250 474854
rect 144486 474618 144528 474854
rect 144208 474586 144528 474618
rect 139088 471454 139408 471486
rect 139088 471218 139130 471454
rect 139366 471218 139408 471454
rect 139088 471134 139408 471218
rect 139088 470898 139130 471134
rect 139366 470898 139408 471134
rect 139088 470866 139408 470898
rect 145794 471454 146414 506898
rect 149328 478894 149648 478926
rect 149328 478658 149370 478894
rect 149606 478658 149648 478894
rect 149328 478574 149648 478658
rect 149328 478338 149370 478574
rect 149606 478338 149648 478574
rect 149328 478306 149648 478338
rect 153234 478894 153854 514338
rect 154448 482614 154768 482646
rect 154448 482378 154490 482614
rect 154726 482378 154768 482614
rect 154448 482294 154768 482378
rect 154448 482058 154490 482294
rect 154726 482058 154768 482294
rect 154448 482026 154768 482058
rect 156954 482614 157574 518058
rect 159568 486334 159888 486366
rect 159568 486098 159610 486334
rect 159846 486098 159888 486334
rect 159568 486014 159888 486098
rect 159568 485778 159610 486014
rect 159846 485778 159888 486014
rect 159568 485746 159888 485778
rect 160674 486334 161294 521778
rect 168114 493774 168734 529218
rect 171834 533494 172454 568938
rect 181794 579454 182414 614898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 602500 186134 618618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 185168 590614 185488 590646
rect 185168 590378 185210 590614
rect 185446 590378 185488 590614
rect 185168 590294 185488 590378
rect 185168 590058 185210 590294
rect 185446 590058 185488 590294
rect 185168 590026 185488 590058
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 180048 550894 180368 550926
rect 180048 550658 180090 550894
rect 180326 550658 180368 550894
rect 180048 550574 180368 550658
rect 180048 550338 180090 550574
rect 180326 550338 180368 550574
rect 180048 550306 180368 550338
rect 174928 547174 175248 547206
rect 174928 546938 174970 547174
rect 175206 546938 175248 547174
rect 174928 546854 175248 546938
rect 174928 546618 174970 546854
rect 175206 546618 175248 546854
rect 174928 546586 175248 546618
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 169808 507454 170128 507486
rect 169808 507218 169850 507454
rect 170086 507218 170128 507454
rect 169808 507134 170128 507218
rect 169808 506898 169850 507134
rect 170086 506898 170128 507134
rect 169808 506866 170128 506898
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 164688 490054 165008 490086
rect 164688 489818 164730 490054
rect 164966 489818 165008 490054
rect 164688 489734 165008 489818
rect 164688 489498 164730 489734
rect 164966 489498 165008 489734
rect 164688 489466 165008 489498
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 133968 454054 134288 454086
rect 133968 453818 134010 454054
rect 134246 453818 134288 454054
rect 133968 453734 134288 453818
rect 133968 453498 134010 453734
rect 134246 453498 134288 453734
rect 133968 453466 134288 453498
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 113488 403174 113808 403206
rect 113488 402938 113530 403174
rect 113766 402938 113808 403174
rect 113488 402854 113808 402938
rect 113488 402618 113530 402854
rect 113766 402618 113808 402854
rect 113488 402586 113808 402618
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 98128 378334 98448 378366
rect 98128 378098 98170 378334
rect 98406 378098 98448 378334
rect 98128 378014 98448 378098
rect 98128 377778 98170 378014
rect 98406 377778 98448 378014
rect 98128 377746 98448 377778
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 93008 338614 93328 338646
rect 93008 338378 93050 338614
rect 93286 338378 93328 338614
rect 93008 338294 93328 338378
rect 93008 338058 93050 338294
rect 93286 338058 93328 338294
rect 93008 338026 93328 338058
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 87888 298894 88208 298926
rect 87888 298658 87930 298894
rect 88166 298658 88208 298894
rect 87888 298574 88208 298658
rect 87888 298338 87930 298574
rect 88166 298338 88208 298574
rect 87888 298306 88208 298338
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 82768 259174 83088 259206
rect 82768 258938 82810 259174
rect 83046 258938 83088 259174
rect 82768 258854 83088 258938
rect 82768 258618 82810 258854
rect 83046 258618 83088 258854
rect 82768 258586 83088 258618
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 72528 202054 72848 202086
rect 72528 201818 72570 202054
rect 72806 201818 72848 202054
rect 72528 201734 72848 201818
rect 72528 201498 72570 201734
rect 72806 201498 72848 201734
rect 72528 201466 72848 201498
rect 67408 198334 67728 198366
rect 67408 198098 67450 198334
rect 67686 198098 67728 198334
rect 67408 198014 67728 198098
rect 67408 197778 67450 198014
rect 67686 197778 67728 198014
rect 67408 197746 67728 197778
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 62288 158614 62608 158646
rect 62288 158378 62330 158614
rect 62566 158378 62608 158614
rect 62288 158294 62608 158378
rect 62288 158058 62330 158294
rect 62566 158058 62608 158294
rect 62288 158026 62608 158058
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 57168 118894 57488 118926
rect 57168 118658 57210 118894
rect 57446 118658 57488 118894
rect 57168 118574 57488 118658
rect 57168 118338 57210 118574
rect 57446 118338 57488 118574
rect 57168 118306 57488 118338
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 56394 58054 57014 93498
rect 60114 97774 60734 133218
rect 63834 137494 64454 172938
rect 73794 183454 74414 218898
rect 77648 219454 77968 219486
rect 77648 219218 77690 219454
rect 77926 219218 77968 219454
rect 77648 219134 77968 219218
rect 77648 218898 77690 219134
rect 77926 218898 77968 219134
rect 77648 218866 77968 218898
rect 81234 190894 81854 226338
rect 84954 230614 85574 266058
rect 88674 270334 89294 305778
rect 96114 313774 96734 349218
rect 99834 353494 100454 388938
rect 103248 382054 103568 382086
rect 103248 381818 103290 382054
rect 103526 381818 103568 382054
rect 103248 381734 103568 381818
rect 103248 381498 103290 381734
rect 103526 381498 103568 381734
rect 103248 381466 103568 381498
rect 108368 363454 108688 363486
rect 108368 363218 108410 363454
rect 108646 363218 108688 363454
rect 108368 363134 108688 363218
rect 108368 362898 108410 363134
rect 108646 362898 108688 363134
rect 108368 362866 108688 362898
rect 109794 363454 110414 398898
rect 117234 370894 117854 406338
rect 118608 406894 118928 406926
rect 118608 406658 118650 406894
rect 118886 406658 118928 406894
rect 118608 406574 118928 406658
rect 118608 406338 118650 406574
rect 118886 406338 118928 406574
rect 118608 406306 118928 406338
rect 120954 374614 121574 410058
rect 123728 410614 124048 410646
rect 123728 410378 123770 410614
rect 124006 410378 124048 410614
rect 123728 410294 124048 410378
rect 123728 410058 123770 410294
rect 124006 410058 124048 410294
rect 123728 410026 124048 410058
rect 124674 378334 125294 413778
rect 128848 414334 129168 414366
rect 128848 414098 128890 414334
rect 129126 414098 129168 414334
rect 128848 414014 129168 414098
rect 128848 413778 128890 414014
rect 129126 413778 129168 414014
rect 128848 413746 129168 413778
rect 132114 385774 132734 421218
rect 135834 425494 136454 460938
rect 144208 439174 144528 439206
rect 144208 438938 144250 439174
rect 144486 438938 144528 439174
rect 144208 438854 144528 438938
rect 144208 438618 144250 438854
rect 144486 438618 144528 438854
rect 144208 438586 144528 438618
rect 139088 435454 139408 435486
rect 139088 435218 139130 435454
rect 139366 435218 139408 435454
rect 139088 435134 139408 435218
rect 139088 434898 139130 435134
rect 139366 434898 139408 435134
rect 139088 434866 139408 434898
rect 145794 435454 146414 470898
rect 149328 442894 149648 442926
rect 149328 442658 149370 442894
rect 149606 442658 149648 442894
rect 149328 442574 149648 442658
rect 149328 442338 149370 442574
rect 149606 442338 149648 442574
rect 149328 442306 149648 442338
rect 153234 442894 153854 478338
rect 154448 446614 154768 446646
rect 154448 446378 154490 446614
rect 154726 446378 154768 446614
rect 154448 446294 154768 446378
rect 154448 446058 154490 446294
rect 154726 446058 154768 446294
rect 154448 446026 154768 446058
rect 156954 446614 157574 482058
rect 159568 450334 159888 450366
rect 159568 450098 159610 450334
rect 159846 450098 159888 450334
rect 159568 450014 159888 450098
rect 159568 449778 159610 450014
rect 159846 449778 159888 450014
rect 159568 449746 159888 449778
rect 160674 450334 161294 485778
rect 168114 457774 168734 493218
rect 171834 497494 172454 532938
rect 181794 543454 182414 578898
rect 189234 586894 189854 622338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 190288 594334 190608 594366
rect 190288 594098 190330 594334
rect 190566 594098 190608 594334
rect 190288 594014 190608 594098
rect 190288 593778 190330 594014
rect 190566 593778 190608 594014
rect 190288 593746 190608 593778
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 185168 554614 185488 554646
rect 185168 554378 185210 554614
rect 185446 554378 185488 554614
rect 185168 554294 185488 554378
rect 185168 554058 185210 554294
rect 185446 554058 185488 554294
rect 185168 554026 185488 554058
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 180048 514894 180368 514926
rect 180048 514658 180090 514894
rect 180326 514658 180368 514894
rect 180048 514574 180368 514658
rect 180048 514338 180090 514574
rect 180326 514338 180368 514574
rect 180048 514306 180368 514338
rect 174928 511174 175248 511206
rect 174928 510938 174970 511174
rect 175206 510938 175248 511174
rect 174928 510854 175248 510938
rect 174928 510618 174970 510854
rect 175206 510618 175248 510854
rect 174928 510586 175248 510618
rect 171834 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 172454 497494
rect 171834 497174 172454 497258
rect 171834 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 172454 497174
rect 169808 471454 170128 471486
rect 169808 471218 169850 471454
rect 170086 471218 170128 471454
rect 169808 471134 170128 471218
rect 169808 470898 169850 471134
rect 170086 470898 170128 471134
rect 169808 470866 170128 470898
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 164688 454054 165008 454086
rect 164688 453818 164730 454054
rect 164966 453818 165008 454054
rect 164688 453734 165008 453818
rect 164688 453498 164730 453734
rect 164966 453498 165008 453734
rect 164688 453466 165008 453498
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 133968 418054 134288 418086
rect 133968 417818 134010 418054
rect 134246 417818 134288 418054
rect 133968 417734 134288 417818
rect 133968 417498 134010 417734
rect 134246 417498 134288 417734
rect 133968 417466 134288 417498
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 113488 367174 113808 367206
rect 113488 366938 113530 367174
rect 113766 366938 113808 367174
rect 113488 366854 113808 366938
rect 113488 366618 113530 366854
rect 113766 366618 113808 366854
rect 113488 366586 113808 366618
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 98128 342334 98448 342366
rect 98128 342098 98170 342334
rect 98406 342098 98448 342334
rect 98128 342014 98448 342098
rect 98128 341778 98170 342014
rect 98406 341778 98448 342014
rect 98128 341746 98448 341778
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 93008 302614 93328 302646
rect 93008 302378 93050 302614
rect 93286 302378 93328 302614
rect 93008 302294 93328 302378
rect 93008 302058 93050 302294
rect 93286 302058 93328 302294
rect 93008 302026 93328 302058
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 87888 262894 88208 262926
rect 87888 262658 87930 262894
rect 88166 262658 88208 262894
rect 87888 262574 88208 262658
rect 87888 262338 87930 262574
rect 88166 262338 88208 262574
rect 87888 262306 88208 262338
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 82768 223174 83088 223206
rect 82768 222938 82810 223174
rect 83046 222938 83088 223174
rect 82768 222854 83088 222938
rect 82768 222618 82810 222854
rect 83046 222618 83088 222854
rect 82768 222586 83088 222618
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 72528 166054 72848 166086
rect 72528 165818 72570 166054
rect 72806 165818 72848 166054
rect 72528 165734 72848 165818
rect 72528 165498 72570 165734
rect 72806 165498 72848 165734
rect 72528 165466 72848 165498
rect 67408 162334 67728 162366
rect 67408 162098 67450 162334
rect 67686 162098 67728 162334
rect 67408 162014 67728 162098
rect 67408 161778 67450 162014
rect 67686 161778 67728 162014
rect 67408 161746 67728 161778
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 62288 122614 62608 122646
rect 62288 122378 62330 122614
rect 62566 122378 62608 122614
rect 62288 122294 62608 122378
rect 62288 122058 62330 122294
rect 62566 122058 62608 122294
rect 62288 122026 62608 122058
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 57168 82894 57488 82926
rect 57168 82658 57210 82894
rect 57446 82658 57488 82894
rect 57168 82574 57488 82658
rect 57168 82338 57210 82574
rect 57446 82338 57488 82574
rect 57168 82306 57488 82338
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 60114 61774 60734 97218
rect 63834 101494 64454 136938
rect 73794 147454 74414 182898
rect 77648 183454 77968 183486
rect 77648 183218 77690 183454
rect 77926 183218 77968 183454
rect 77648 183134 77968 183218
rect 77648 182898 77690 183134
rect 77926 182898 77968 183134
rect 77648 182866 77968 182898
rect 81234 154894 81854 190338
rect 84954 194614 85574 230058
rect 88674 234334 89294 269778
rect 96114 277774 96734 313218
rect 99834 317494 100454 352938
rect 103248 346054 103568 346086
rect 103248 345818 103290 346054
rect 103526 345818 103568 346054
rect 103248 345734 103568 345818
rect 103248 345498 103290 345734
rect 103526 345498 103568 345734
rect 103248 345466 103568 345498
rect 108368 327454 108688 327486
rect 108368 327218 108410 327454
rect 108646 327218 108688 327454
rect 108368 327134 108688 327218
rect 108368 326898 108410 327134
rect 108646 326898 108688 327134
rect 108368 326866 108688 326898
rect 109794 327454 110414 362898
rect 117234 334894 117854 370338
rect 118608 370894 118928 370926
rect 118608 370658 118650 370894
rect 118886 370658 118928 370894
rect 118608 370574 118928 370658
rect 118608 370338 118650 370574
rect 118886 370338 118928 370574
rect 118608 370306 118928 370338
rect 120954 338614 121574 374058
rect 123728 374614 124048 374646
rect 123728 374378 123770 374614
rect 124006 374378 124048 374614
rect 123728 374294 124048 374378
rect 123728 374058 123770 374294
rect 124006 374058 124048 374294
rect 123728 374026 124048 374058
rect 124674 342334 125294 377778
rect 128848 378334 129168 378366
rect 128848 378098 128890 378334
rect 129126 378098 129168 378334
rect 128848 378014 129168 378098
rect 128848 377778 128890 378014
rect 129126 377778 129168 378014
rect 128848 377746 129168 377778
rect 132114 349774 132734 385218
rect 135834 389494 136454 424938
rect 144208 403174 144528 403206
rect 144208 402938 144250 403174
rect 144486 402938 144528 403174
rect 144208 402854 144528 402938
rect 144208 402618 144250 402854
rect 144486 402618 144528 402854
rect 144208 402586 144528 402618
rect 139088 399454 139408 399486
rect 139088 399218 139130 399454
rect 139366 399218 139408 399454
rect 139088 399134 139408 399218
rect 139088 398898 139130 399134
rect 139366 398898 139408 399134
rect 139088 398866 139408 398898
rect 145794 399454 146414 434898
rect 149328 406894 149648 406926
rect 149328 406658 149370 406894
rect 149606 406658 149648 406894
rect 149328 406574 149648 406658
rect 149328 406338 149370 406574
rect 149606 406338 149648 406574
rect 149328 406306 149648 406338
rect 153234 406894 153854 442338
rect 154448 410614 154768 410646
rect 154448 410378 154490 410614
rect 154726 410378 154768 410614
rect 154448 410294 154768 410378
rect 154448 410058 154490 410294
rect 154726 410058 154768 410294
rect 154448 410026 154768 410058
rect 156954 410614 157574 446058
rect 159568 414334 159888 414366
rect 159568 414098 159610 414334
rect 159846 414098 159888 414334
rect 159568 414014 159888 414098
rect 159568 413778 159610 414014
rect 159846 413778 159888 414014
rect 159568 413746 159888 413778
rect 160674 414334 161294 449778
rect 168114 421774 168734 457218
rect 171834 461494 172454 496938
rect 181794 507454 182414 542898
rect 189234 550894 189854 586338
rect 192954 590614 193574 626058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 195408 598054 195728 598086
rect 195408 597818 195450 598054
rect 195686 597818 195728 598054
rect 195408 597734 195728 597818
rect 195408 597498 195450 597734
rect 195686 597498 195728 597734
rect 195408 597466 195728 597498
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 190288 558334 190608 558366
rect 190288 558098 190330 558334
rect 190566 558098 190608 558334
rect 190288 558014 190608 558098
rect 190288 557778 190330 558014
rect 190566 557778 190608 558014
rect 190288 557746 190608 557778
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 185168 518614 185488 518646
rect 185168 518378 185210 518614
rect 185446 518378 185488 518614
rect 185168 518294 185488 518378
rect 185168 518058 185210 518294
rect 185446 518058 185488 518294
rect 185168 518026 185488 518058
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 180048 478894 180368 478926
rect 180048 478658 180090 478894
rect 180326 478658 180368 478894
rect 180048 478574 180368 478658
rect 180048 478338 180090 478574
rect 180326 478338 180368 478574
rect 180048 478306 180368 478338
rect 174928 475174 175248 475206
rect 174928 474938 174970 475174
rect 175206 474938 175248 475174
rect 174928 474854 175248 474938
rect 174928 474618 174970 474854
rect 175206 474618 175248 474854
rect 174928 474586 175248 474618
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 169808 435454 170128 435486
rect 169808 435218 169850 435454
rect 170086 435218 170128 435454
rect 169808 435134 170128 435218
rect 169808 434898 169850 435134
rect 170086 434898 170128 435134
rect 169808 434866 170128 434898
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 164688 418054 165008 418086
rect 164688 417818 164730 418054
rect 164966 417818 165008 418054
rect 164688 417734 165008 417818
rect 164688 417498 164730 417734
rect 164966 417498 165008 417734
rect 164688 417466 165008 417498
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 133968 382054 134288 382086
rect 133968 381818 134010 382054
rect 134246 381818 134288 382054
rect 133968 381734 134288 381818
rect 133968 381498 134010 381734
rect 134246 381498 134288 381734
rect 133968 381466 134288 381498
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 113488 331174 113808 331206
rect 113488 330938 113530 331174
rect 113766 330938 113808 331174
rect 113488 330854 113808 330938
rect 113488 330618 113530 330854
rect 113766 330618 113808 330854
rect 113488 330586 113808 330618
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 98128 306334 98448 306366
rect 98128 306098 98170 306334
rect 98406 306098 98448 306334
rect 98128 306014 98448 306098
rect 98128 305778 98170 306014
rect 98406 305778 98448 306014
rect 98128 305746 98448 305778
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 93008 266614 93328 266646
rect 93008 266378 93050 266614
rect 93286 266378 93328 266614
rect 93008 266294 93328 266378
rect 93008 266058 93050 266294
rect 93286 266058 93328 266294
rect 93008 266026 93328 266058
rect 88674 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 89294 234334
rect 88674 234014 89294 234098
rect 88674 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 89294 234014
rect 87888 226894 88208 226926
rect 87888 226658 87930 226894
rect 88166 226658 88208 226894
rect 87888 226574 88208 226658
rect 87888 226338 87930 226574
rect 88166 226338 88208 226574
rect 87888 226306 88208 226338
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 82768 187174 83088 187206
rect 82768 186938 82810 187174
rect 83046 186938 83088 187174
rect 82768 186854 83088 186938
rect 82768 186618 82810 186854
rect 83046 186618 83088 186854
rect 82768 186586 83088 186618
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 72528 130054 72848 130086
rect 72528 129818 72570 130054
rect 72806 129818 72848 130054
rect 72528 129734 72848 129818
rect 72528 129498 72570 129734
rect 72806 129498 72848 129734
rect 72528 129466 72848 129498
rect 67408 126334 67728 126366
rect 67408 126098 67450 126334
rect 67686 126098 67728 126334
rect 67408 126014 67728 126098
rect 67408 125778 67450 126014
rect 67686 125778 67728 126014
rect 67408 125746 67728 125778
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 62288 86614 62608 86646
rect 62288 86378 62330 86614
rect 62566 86378 62608 86614
rect 62288 86294 62608 86378
rect 62288 86058 62330 86294
rect 62566 86058 62608 86294
rect 62288 86026 62608 86058
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 57168 46894 57488 46926
rect 57168 46658 57210 46894
rect 57446 46658 57488 46894
rect 57168 46574 57488 46658
rect 57168 46338 57210 46574
rect 57446 46338 57488 46574
rect 57168 46306 57488 46338
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 60114 25774 60734 61218
rect 63834 65494 64454 100938
rect 73794 111454 74414 146898
rect 77648 147454 77968 147486
rect 77648 147218 77690 147454
rect 77926 147218 77968 147454
rect 77648 147134 77968 147218
rect 77648 146898 77690 147134
rect 77926 146898 77968 147134
rect 77648 146866 77968 146898
rect 81234 118894 81854 154338
rect 84954 158614 85574 194058
rect 88674 198334 89294 233778
rect 96114 241774 96734 277218
rect 99834 281494 100454 316938
rect 103248 310054 103568 310086
rect 103248 309818 103290 310054
rect 103526 309818 103568 310054
rect 103248 309734 103568 309818
rect 103248 309498 103290 309734
rect 103526 309498 103568 309734
rect 103248 309466 103568 309498
rect 108368 291454 108688 291486
rect 108368 291218 108410 291454
rect 108646 291218 108688 291454
rect 108368 291134 108688 291218
rect 108368 290898 108410 291134
rect 108646 290898 108688 291134
rect 108368 290866 108688 290898
rect 109794 291454 110414 326898
rect 117234 298894 117854 334338
rect 118608 334894 118928 334926
rect 118608 334658 118650 334894
rect 118886 334658 118928 334894
rect 118608 334574 118928 334658
rect 118608 334338 118650 334574
rect 118886 334338 118928 334574
rect 118608 334306 118928 334338
rect 120954 302614 121574 338058
rect 123728 338614 124048 338646
rect 123728 338378 123770 338614
rect 124006 338378 124048 338614
rect 123728 338294 124048 338378
rect 123728 338058 123770 338294
rect 124006 338058 124048 338294
rect 123728 338026 124048 338058
rect 124674 306334 125294 341778
rect 128848 342334 129168 342366
rect 128848 342098 128890 342334
rect 129126 342098 129168 342334
rect 128848 342014 129168 342098
rect 128848 341778 128890 342014
rect 129126 341778 129168 342014
rect 128848 341746 129168 341778
rect 132114 313774 132734 349218
rect 135834 353494 136454 388938
rect 144208 367174 144528 367206
rect 144208 366938 144250 367174
rect 144486 366938 144528 367174
rect 144208 366854 144528 366938
rect 144208 366618 144250 366854
rect 144486 366618 144528 366854
rect 144208 366586 144528 366618
rect 139088 363454 139408 363486
rect 139088 363218 139130 363454
rect 139366 363218 139408 363454
rect 139088 363134 139408 363218
rect 139088 362898 139130 363134
rect 139366 362898 139408 363134
rect 139088 362866 139408 362898
rect 145794 363454 146414 398898
rect 149328 370894 149648 370926
rect 149328 370658 149370 370894
rect 149606 370658 149648 370894
rect 149328 370574 149648 370658
rect 149328 370338 149370 370574
rect 149606 370338 149648 370574
rect 149328 370306 149648 370338
rect 153234 370894 153854 406338
rect 154448 374614 154768 374646
rect 154448 374378 154490 374614
rect 154726 374378 154768 374614
rect 154448 374294 154768 374378
rect 154448 374058 154490 374294
rect 154726 374058 154768 374294
rect 154448 374026 154768 374058
rect 156954 374614 157574 410058
rect 159568 378334 159888 378366
rect 159568 378098 159610 378334
rect 159846 378098 159888 378334
rect 159568 378014 159888 378098
rect 159568 377778 159610 378014
rect 159846 377778 159888 378014
rect 159568 377746 159888 377778
rect 160674 378334 161294 413778
rect 168114 385774 168734 421218
rect 171834 425494 172454 460938
rect 181794 471454 182414 506898
rect 189234 514894 189854 550338
rect 192954 554614 193574 590058
rect 196674 594334 197294 629778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 602500 201014 633498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 195408 562054 195728 562086
rect 195408 561818 195450 562054
rect 195686 561818 195728 562054
rect 195408 561734 195728 561818
rect 195408 561498 195450 561734
rect 195686 561498 195728 561734
rect 195408 561466 195728 561498
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 190288 522334 190608 522366
rect 190288 522098 190330 522334
rect 190566 522098 190608 522334
rect 190288 522014 190608 522098
rect 190288 521778 190330 522014
rect 190566 521778 190608 522014
rect 190288 521746 190608 521778
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 185168 482614 185488 482646
rect 185168 482378 185210 482614
rect 185446 482378 185488 482614
rect 185168 482294 185488 482378
rect 185168 482058 185210 482294
rect 185446 482058 185488 482294
rect 185168 482026 185488 482058
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 180048 442894 180368 442926
rect 180048 442658 180090 442894
rect 180326 442658 180368 442894
rect 180048 442574 180368 442658
rect 180048 442338 180090 442574
rect 180326 442338 180368 442574
rect 180048 442306 180368 442338
rect 174928 439174 175248 439206
rect 174928 438938 174970 439174
rect 175206 438938 175248 439174
rect 174928 438854 175248 438938
rect 174928 438618 174970 438854
rect 175206 438618 175248 438854
rect 174928 438586 175248 438618
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 169808 399454 170128 399486
rect 169808 399218 169850 399454
rect 170086 399218 170128 399454
rect 169808 399134 170128 399218
rect 169808 398898 169850 399134
rect 170086 398898 170128 399134
rect 169808 398866 170128 398898
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 164688 382054 165008 382086
rect 164688 381818 164730 382054
rect 164966 381818 165008 382054
rect 164688 381734 165008 381818
rect 164688 381498 164730 381734
rect 164966 381498 165008 381734
rect 164688 381466 165008 381498
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 133968 346054 134288 346086
rect 133968 345818 134010 346054
rect 134246 345818 134288 346054
rect 133968 345734 134288 345818
rect 133968 345498 134010 345734
rect 134246 345498 134288 345734
rect 133968 345466 134288 345498
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 113488 295174 113808 295206
rect 113488 294938 113530 295174
rect 113766 294938 113808 295174
rect 113488 294854 113808 294938
rect 113488 294618 113530 294854
rect 113766 294618 113808 294854
rect 113488 294586 113808 294618
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 99834 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 100454 281494
rect 99834 281174 100454 281258
rect 99834 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 100454 281174
rect 98128 270334 98448 270366
rect 98128 270098 98170 270334
rect 98406 270098 98448 270334
rect 98128 270014 98448 270098
rect 98128 269778 98170 270014
rect 98406 269778 98448 270014
rect 98128 269746 98448 269778
rect 96114 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 96734 241774
rect 96114 241454 96734 241538
rect 96114 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 96734 241454
rect 93008 230614 93328 230646
rect 93008 230378 93050 230614
rect 93286 230378 93328 230614
rect 93008 230294 93328 230378
rect 93008 230058 93050 230294
rect 93286 230058 93328 230294
rect 93008 230026 93328 230058
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 87888 190894 88208 190926
rect 87888 190658 87930 190894
rect 88166 190658 88208 190894
rect 87888 190574 88208 190658
rect 87888 190338 87930 190574
rect 88166 190338 88208 190574
rect 87888 190306 88208 190338
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 82768 151174 83088 151206
rect 82768 150938 82810 151174
rect 83046 150938 83088 151174
rect 82768 150854 83088 150938
rect 82768 150618 82810 150854
rect 83046 150618 83088 150854
rect 82768 150586 83088 150618
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 72528 94054 72848 94086
rect 72528 93818 72570 94054
rect 72806 93818 72848 94054
rect 72528 93734 72848 93818
rect 72528 93498 72570 93734
rect 72806 93498 72848 93734
rect 72528 93466 72848 93498
rect 67408 90334 67728 90366
rect 67408 90098 67450 90334
rect 67686 90098 67728 90334
rect 67408 90014 67728 90098
rect 67408 89778 67450 90014
rect 67686 89778 67728 90014
rect 67408 89746 67728 89778
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 62288 50614 62608 50646
rect 62288 50378 62330 50614
rect 62566 50378 62608 50614
rect 62288 50294 62608 50378
rect 62288 50058 62330 50294
rect 62566 50058 62608 50294
rect 62288 50026 62608 50058
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 57168 10894 57488 10926
rect 57168 10658 57210 10894
rect 57446 10658 57488 10894
rect 57168 10574 57488 10658
rect 57168 10338 57210 10574
rect 57446 10338 57488 10574
rect 57168 10306 57488 10338
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 -6106 60734 25218
rect 63834 29494 64454 64938
rect 73794 75454 74414 110898
rect 77648 111454 77968 111486
rect 77648 111218 77690 111454
rect 77926 111218 77968 111454
rect 77648 111134 77968 111218
rect 77648 110898 77690 111134
rect 77926 110898 77968 111134
rect 77648 110866 77968 110898
rect 81234 82894 81854 118338
rect 84954 122614 85574 158058
rect 88674 162334 89294 197778
rect 96114 205774 96734 241218
rect 99834 245494 100454 280938
rect 103248 274054 103568 274086
rect 103248 273818 103290 274054
rect 103526 273818 103568 274054
rect 103248 273734 103568 273818
rect 103248 273498 103290 273734
rect 103526 273498 103568 273734
rect 103248 273466 103568 273498
rect 108368 255454 108688 255486
rect 108368 255218 108410 255454
rect 108646 255218 108688 255454
rect 108368 255134 108688 255218
rect 108368 254898 108410 255134
rect 108646 254898 108688 255134
rect 108368 254866 108688 254898
rect 109794 255454 110414 290898
rect 117234 262894 117854 298338
rect 118608 298894 118928 298926
rect 118608 298658 118650 298894
rect 118886 298658 118928 298894
rect 118608 298574 118928 298658
rect 118608 298338 118650 298574
rect 118886 298338 118928 298574
rect 118608 298306 118928 298338
rect 120954 266614 121574 302058
rect 123728 302614 124048 302646
rect 123728 302378 123770 302614
rect 124006 302378 124048 302614
rect 123728 302294 124048 302378
rect 123728 302058 123770 302294
rect 124006 302058 124048 302294
rect 123728 302026 124048 302058
rect 124674 270334 125294 305778
rect 128848 306334 129168 306366
rect 128848 306098 128890 306334
rect 129126 306098 129168 306334
rect 128848 306014 129168 306098
rect 128848 305778 128890 306014
rect 129126 305778 129168 306014
rect 128848 305746 129168 305778
rect 132114 277774 132734 313218
rect 135834 317494 136454 352938
rect 144208 331174 144528 331206
rect 144208 330938 144250 331174
rect 144486 330938 144528 331174
rect 144208 330854 144528 330938
rect 144208 330618 144250 330854
rect 144486 330618 144528 330854
rect 144208 330586 144528 330618
rect 139088 327454 139408 327486
rect 139088 327218 139130 327454
rect 139366 327218 139408 327454
rect 139088 327134 139408 327218
rect 139088 326898 139130 327134
rect 139366 326898 139408 327134
rect 139088 326866 139408 326898
rect 145794 327454 146414 362898
rect 149328 334894 149648 334926
rect 149328 334658 149370 334894
rect 149606 334658 149648 334894
rect 149328 334574 149648 334658
rect 149328 334338 149370 334574
rect 149606 334338 149648 334574
rect 149328 334306 149648 334338
rect 153234 334894 153854 370338
rect 154448 338614 154768 338646
rect 154448 338378 154490 338614
rect 154726 338378 154768 338614
rect 154448 338294 154768 338378
rect 154448 338058 154490 338294
rect 154726 338058 154768 338294
rect 154448 338026 154768 338058
rect 156954 338614 157574 374058
rect 159568 342334 159888 342366
rect 159568 342098 159610 342334
rect 159846 342098 159888 342334
rect 159568 342014 159888 342098
rect 159568 341778 159610 342014
rect 159846 341778 159888 342014
rect 159568 341746 159888 341778
rect 160674 342334 161294 377778
rect 168114 349774 168734 385218
rect 171834 389494 172454 424938
rect 181794 435454 182414 470898
rect 189234 478894 189854 514338
rect 192954 518614 193574 554058
rect 196674 558334 197294 593778
rect 204114 601774 204734 637218
rect 204114 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 204734 601774
rect 204114 601454 204734 601538
rect 204114 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 204734 601454
rect 200528 579454 200848 579486
rect 200528 579218 200570 579454
rect 200806 579218 200848 579454
rect 200528 579134 200848 579218
rect 200528 578898 200570 579134
rect 200806 578898 200848 579134
rect 200528 578866 200848 578898
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 195408 526054 195728 526086
rect 195408 525818 195450 526054
rect 195686 525818 195728 526054
rect 195408 525734 195728 525818
rect 195408 525498 195450 525734
rect 195686 525498 195728 525734
rect 195408 525466 195728 525498
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 190288 486334 190608 486366
rect 190288 486098 190330 486334
rect 190566 486098 190608 486334
rect 190288 486014 190608 486098
rect 190288 485778 190330 486014
rect 190566 485778 190608 486014
rect 190288 485746 190608 485778
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 185168 446614 185488 446646
rect 185168 446378 185210 446614
rect 185446 446378 185488 446614
rect 185168 446294 185488 446378
rect 185168 446058 185210 446294
rect 185446 446058 185488 446294
rect 185168 446026 185488 446058
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 180048 406894 180368 406926
rect 180048 406658 180090 406894
rect 180326 406658 180368 406894
rect 180048 406574 180368 406658
rect 180048 406338 180090 406574
rect 180326 406338 180368 406574
rect 180048 406306 180368 406338
rect 174928 403174 175248 403206
rect 174928 402938 174970 403174
rect 175206 402938 175248 403174
rect 174928 402854 175248 402938
rect 174928 402618 174970 402854
rect 175206 402618 175248 402854
rect 174928 402586 175248 402618
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 169808 363454 170128 363486
rect 169808 363218 169850 363454
rect 170086 363218 170128 363454
rect 169808 363134 170128 363218
rect 169808 362898 169850 363134
rect 170086 362898 170128 363134
rect 169808 362866 170128 362898
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 164688 346054 165008 346086
rect 164688 345818 164730 346054
rect 164966 345818 165008 346054
rect 164688 345734 165008 345818
rect 164688 345498 164730 345734
rect 164966 345498 165008 345734
rect 164688 345466 165008 345498
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 133968 310054 134288 310086
rect 133968 309818 134010 310054
rect 134246 309818 134288 310054
rect 133968 309734 134288 309818
rect 133968 309498 134010 309734
rect 134246 309498 134288 309734
rect 133968 309466 134288 309498
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 113488 259174 113808 259206
rect 113488 258938 113530 259174
rect 113766 258938 113808 259174
rect 113488 258854 113808 258938
rect 113488 258618 113530 258854
rect 113766 258618 113808 258854
rect 113488 258586 113808 258618
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 99834 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 100454 245494
rect 99834 245174 100454 245258
rect 99834 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 100454 245174
rect 98128 234334 98448 234366
rect 98128 234098 98170 234334
rect 98406 234098 98448 234334
rect 98128 234014 98448 234098
rect 98128 233778 98170 234014
rect 98406 233778 98448 234014
rect 98128 233746 98448 233778
rect 96114 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 96734 205774
rect 96114 205454 96734 205538
rect 96114 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 96734 205454
rect 93008 194614 93328 194646
rect 93008 194378 93050 194614
rect 93286 194378 93328 194614
rect 93008 194294 93328 194378
rect 93008 194058 93050 194294
rect 93286 194058 93328 194294
rect 93008 194026 93328 194058
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 87888 154894 88208 154926
rect 87888 154658 87930 154894
rect 88166 154658 88208 154894
rect 87888 154574 88208 154658
rect 87888 154338 87930 154574
rect 88166 154338 88208 154574
rect 87888 154306 88208 154338
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 82768 115174 83088 115206
rect 82768 114938 82810 115174
rect 83046 114938 83088 115174
rect 82768 114854 83088 114938
rect 82768 114618 82810 114854
rect 83046 114618 83088 114854
rect 82768 114586 83088 114618
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 72528 58054 72848 58086
rect 72528 57818 72570 58054
rect 72806 57818 72848 58054
rect 72528 57734 72848 57818
rect 72528 57498 72570 57734
rect 72806 57498 72848 57734
rect 72528 57466 72848 57498
rect 67408 54334 67728 54366
rect 67408 54098 67450 54334
rect 67686 54098 67728 54334
rect 67408 54014 67728 54098
rect 67408 53778 67450 54014
rect 67686 53778 67728 54014
rect 67408 53746 67728 53778
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 62288 14614 62608 14646
rect 62288 14378 62330 14614
rect 62566 14378 62608 14614
rect 62288 14294 62608 14378
rect 62288 14058 62330 14294
rect 62566 14058 62608 14294
rect 62288 14026 62608 14058
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 -7066 64454 28938
rect 73794 39454 74414 74898
rect 77648 75454 77968 75486
rect 77648 75218 77690 75454
rect 77926 75218 77968 75454
rect 77648 75134 77968 75218
rect 77648 74898 77690 75134
rect 77926 74898 77968 75134
rect 77648 74866 77968 74898
rect 81234 46894 81854 82338
rect 84954 86614 85574 122058
rect 88674 126334 89294 161778
rect 96114 169774 96734 205218
rect 99834 209494 100454 244938
rect 103248 238054 103568 238086
rect 103248 237818 103290 238054
rect 103526 237818 103568 238054
rect 103248 237734 103568 237818
rect 103248 237498 103290 237734
rect 103526 237498 103568 237734
rect 103248 237466 103568 237498
rect 108368 219454 108688 219486
rect 108368 219218 108410 219454
rect 108646 219218 108688 219454
rect 108368 219134 108688 219218
rect 108368 218898 108410 219134
rect 108646 218898 108688 219134
rect 108368 218866 108688 218898
rect 109794 219454 110414 254898
rect 117234 226894 117854 262338
rect 118608 262894 118928 262926
rect 118608 262658 118650 262894
rect 118886 262658 118928 262894
rect 118608 262574 118928 262658
rect 118608 262338 118650 262574
rect 118886 262338 118928 262574
rect 118608 262306 118928 262338
rect 120954 230614 121574 266058
rect 123728 266614 124048 266646
rect 123728 266378 123770 266614
rect 124006 266378 124048 266614
rect 123728 266294 124048 266378
rect 123728 266058 123770 266294
rect 124006 266058 124048 266294
rect 123728 266026 124048 266058
rect 124674 234334 125294 269778
rect 128848 270334 129168 270366
rect 128848 270098 128890 270334
rect 129126 270098 129168 270334
rect 128848 270014 129168 270098
rect 128848 269778 128890 270014
rect 129126 269778 129168 270014
rect 128848 269746 129168 269778
rect 132114 241774 132734 277218
rect 135834 281494 136454 316938
rect 144208 295174 144528 295206
rect 144208 294938 144250 295174
rect 144486 294938 144528 295174
rect 144208 294854 144528 294938
rect 144208 294618 144250 294854
rect 144486 294618 144528 294854
rect 144208 294586 144528 294618
rect 139088 291454 139408 291486
rect 139088 291218 139130 291454
rect 139366 291218 139408 291454
rect 139088 291134 139408 291218
rect 139088 290898 139130 291134
rect 139366 290898 139408 291134
rect 139088 290866 139408 290898
rect 145794 291454 146414 326898
rect 149328 298894 149648 298926
rect 149328 298658 149370 298894
rect 149606 298658 149648 298894
rect 149328 298574 149648 298658
rect 149328 298338 149370 298574
rect 149606 298338 149648 298574
rect 149328 298306 149648 298338
rect 153234 298894 153854 334338
rect 154448 302614 154768 302646
rect 154448 302378 154490 302614
rect 154726 302378 154768 302614
rect 154448 302294 154768 302378
rect 154448 302058 154490 302294
rect 154726 302058 154768 302294
rect 154448 302026 154768 302058
rect 156954 302614 157574 338058
rect 159568 306334 159888 306366
rect 159568 306098 159610 306334
rect 159846 306098 159888 306334
rect 159568 306014 159888 306098
rect 159568 305778 159610 306014
rect 159846 305778 159888 306014
rect 159568 305746 159888 305778
rect 160674 306334 161294 341778
rect 168114 313774 168734 349218
rect 171834 353494 172454 388938
rect 181794 399454 182414 434898
rect 189234 442894 189854 478338
rect 192954 482614 193574 518058
rect 196674 522334 197294 557778
rect 204114 565774 204734 601218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 205648 583174 205968 583206
rect 205648 582938 205690 583174
rect 205926 582938 205968 583174
rect 205648 582854 205968 582938
rect 205648 582618 205690 582854
rect 205926 582618 205968 582854
rect 205648 582586 205968 582618
rect 204114 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 204734 565774
rect 204114 565454 204734 565538
rect 204114 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 204734 565454
rect 200528 543454 200848 543486
rect 200528 543218 200570 543454
rect 200806 543218 200848 543454
rect 200528 543134 200848 543218
rect 200528 542898 200570 543134
rect 200806 542898 200848 543134
rect 200528 542866 200848 542898
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 195408 490054 195728 490086
rect 195408 489818 195450 490054
rect 195686 489818 195728 490054
rect 195408 489734 195728 489818
rect 195408 489498 195450 489734
rect 195686 489498 195728 489734
rect 195408 489466 195728 489498
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190288 450334 190608 450366
rect 190288 450098 190330 450334
rect 190566 450098 190608 450334
rect 190288 450014 190608 450098
rect 190288 449778 190330 450014
rect 190566 449778 190608 450014
rect 190288 449746 190608 449778
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 185168 410614 185488 410646
rect 185168 410378 185210 410614
rect 185446 410378 185488 410614
rect 185168 410294 185488 410378
rect 185168 410058 185210 410294
rect 185446 410058 185488 410294
rect 185168 410026 185488 410058
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 180048 370894 180368 370926
rect 180048 370658 180090 370894
rect 180326 370658 180368 370894
rect 180048 370574 180368 370658
rect 180048 370338 180090 370574
rect 180326 370338 180368 370574
rect 180048 370306 180368 370338
rect 174928 367174 175248 367206
rect 174928 366938 174970 367174
rect 175206 366938 175248 367174
rect 174928 366854 175248 366938
rect 174928 366618 174970 366854
rect 175206 366618 175248 366854
rect 174928 366586 175248 366618
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 169808 327454 170128 327486
rect 169808 327218 169850 327454
rect 170086 327218 170128 327454
rect 169808 327134 170128 327218
rect 169808 326898 169850 327134
rect 170086 326898 170128 327134
rect 169808 326866 170128 326898
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 164688 310054 165008 310086
rect 164688 309818 164730 310054
rect 164966 309818 165008 310054
rect 164688 309734 165008 309818
rect 164688 309498 164730 309734
rect 164966 309498 165008 309734
rect 164688 309466 165008 309498
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 133968 274054 134288 274086
rect 133968 273818 134010 274054
rect 134246 273818 134288 274054
rect 133968 273734 134288 273818
rect 133968 273498 134010 273734
rect 134246 273498 134288 273734
rect 133968 273466 134288 273498
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 113488 223174 113808 223206
rect 113488 222938 113530 223174
rect 113766 222938 113808 223174
rect 113488 222854 113808 222938
rect 113488 222618 113530 222854
rect 113766 222618 113808 222854
rect 113488 222586 113808 222618
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 99834 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 100454 209494
rect 99834 209174 100454 209258
rect 99834 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 100454 209174
rect 98128 198334 98448 198366
rect 98128 198098 98170 198334
rect 98406 198098 98448 198334
rect 98128 198014 98448 198098
rect 98128 197778 98170 198014
rect 98406 197778 98448 198014
rect 98128 197746 98448 197778
rect 96114 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 96734 169774
rect 96114 169454 96734 169538
rect 96114 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 96734 169454
rect 93008 158614 93328 158646
rect 93008 158378 93050 158614
rect 93286 158378 93328 158614
rect 93008 158294 93328 158378
rect 93008 158058 93050 158294
rect 93286 158058 93328 158294
rect 93008 158026 93328 158058
rect 88674 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 89294 126334
rect 88674 126014 89294 126098
rect 88674 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 89294 126014
rect 87888 118894 88208 118926
rect 87888 118658 87930 118894
rect 88166 118658 88208 118894
rect 87888 118574 88208 118658
rect 87888 118338 87930 118574
rect 88166 118338 88208 118574
rect 87888 118306 88208 118338
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 82768 79174 83088 79206
rect 82768 78938 82810 79174
rect 83046 78938 83088 79174
rect 82768 78854 83088 78938
rect 82768 78618 82810 78854
rect 83046 78618 83088 78854
rect 82768 78586 83088 78618
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 72528 22054 72848 22086
rect 72528 21818 72570 22054
rect 72806 21818 72848 22054
rect 72528 21734 72848 21818
rect 72528 21498 72570 21734
rect 72806 21498 72848 21734
rect 72528 21466 72848 21498
rect 67408 18334 67728 18366
rect 67408 18098 67450 18334
rect 67686 18098 67728 18334
rect 67408 18014 67728 18098
rect 67408 17778 67450 18014
rect 67686 17778 67728 18014
rect 67408 17746 67728 17778
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 3454 74414 38898
rect 77648 39454 77968 39486
rect 77648 39218 77690 39454
rect 77926 39218 77968 39454
rect 77648 39134 77968 39218
rect 77648 38898 77690 39134
rect 77926 38898 77968 39134
rect 77648 38866 77968 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 81234 10894 81854 46338
rect 84954 50614 85574 86058
rect 88674 90334 89294 125778
rect 96114 133774 96734 169218
rect 99834 173494 100454 208938
rect 103248 202054 103568 202086
rect 103248 201818 103290 202054
rect 103526 201818 103568 202054
rect 103248 201734 103568 201818
rect 103248 201498 103290 201734
rect 103526 201498 103568 201734
rect 103248 201466 103568 201498
rect 108368 183454 108688 183486
rect 108368 183218 108410 183454
rect 108646 183218 108688 183454
rect 108368 183134 108688 183218
rect 108368 182898 108410 183134
rect 108646 182898 108688 183134
rect 108368 182866 108688 182898
rect 109794 183454 110414 218898
rect 117234 190894 117854 226338
rect 118608 226894 118928 226926
rect 118608 226658 118650 226894
rect 118886 226658 118928 226894
rect 118608 226574 118928 226658
rect 118608 226338 118650 226574
rect 118886 226338 118928 226574
rect 118608 226306 118928 226338
rect 120954 194614 121574 230058
rect 123728 230614 124048 230646
rect 123728 230378 123770 230614
rect 124006 230378 124048 230614
rect 123728 230294 124048 230378
rect 123728 230058 123770 230294
rect 124006 230058 124048 230294
rect 123728 230026 124048 230058
rect 124674 198334 125294 233778
rect 128848 234334 129168 234366
rect 128848 234098 128890 234334
rect 129126 234098 129168 234334
rect 128848 234014 129168 234098
rect 128848 233778 128890 234014
rect 129126 233778 129168 234014
rect 128848 233746 129168 233778
rect 132114 205774 132734 241218
rect 135834 245494 136454 280938
rect 144208 259174 144528 259206
rect 144208 258938 144250 259174
rect 144486 258938 144528 259174
rect 144208 258854 144528 258938
rect 144208 258618 144250 258854
rect 144486 258618 144528 258854
rect 144208 258586 144528 258618
rect 139088 255454 139408 255486
rect 139088 255218 139130 255454
rect 139366 255218 139408 255454
rect 139088 255134 139408 255218
rect 139088 254898 139130 255134
rect 139366 254898 139408 255134
rect 139088 254866 139408 254898
rect 145794 255454 146414 290898
rect 149328 262894 149648 262926
rect 149328 262658 149370 262894
rect 149606 262658 149648 262894
rect 149328 262574 149648 262658
rect 149328 262338 149370 262574
rect 149606 262338 149648 262574
rect 149328 262306 149648 262338
rect 153234 262894 153854 298338
rect 154448 266614 154768 266646
rect 154448 266378 154490 266614
rect 154726 266378 154768 266614
rect 154448 266294 154768 266378
rect 154448 266058 154490 266294
rect 154726 266058 154768 266294
rect 154448 266026 154768 266058
rect 156954 266614 157574 302058
rect 159568 270334 159888 270366
rect 159568 270098 159610 270334
rect 159846 270098 159888 270334
rect 159568 270014 159888 270098
rect 159568 269778 159610 270014
rect 159846 269778 159888 270014
rect 159568 269746 159888 269778
rect 160674 270334 161294 305778
rect 168114 277774 168734 313218
rect 171834 317494 172454 352938
rect 181794 363454 182414 398898
rect 189234 406894 189854 442338
rect 192954 446614 193574 482058
rect 196674 486334 197294 521778
rect 204114 529774 204734 565218
rect 207834 569494 208454 604938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 215888 590614 216208 590646
rect 215888 590378 215930 590614
rect 216166 590378 216208 590614
rect 215888 590294 216208 590378
rect 215888 590058 215930 590294
rect 216166 590058 216208 590294
rect 215888 590026 216208 590058
rect 210768 586894 211088 586926
rect 210768 586658 210810 586894
rect 211046 586658 211088 586894
rect 210768 586574 211088 586658
rect 210768 586338 210810 586574
rect 211046 586338 211088 586574
rect 210768 586306 211088 586338
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 205648 547174 205968 547206
rect 205648 546938 205690 547174
rect 205926 546938 205968 547174
rect 205648 546854 205968 546938
rect 205648 546618 205690 546854
rect 205926 546618 205968 546854
rect 205648 546586 205968 546618
rect 204114 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 204734 529774
rect 204114 529454 204734 529538
rect 204114 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 204734 529454
rect 200528 507454 200848 507486
rect 200528 507218 200570 507454
rect 200806 507218 200848 507454
rect 200528 507134 200848 507218
rect 200528 506898 200570 507134
rect 200806 506898 200848 507134
rect 200528 506866 200848 506898
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 195408 454054 195728 454086
rect 195408 453818 195450 454054
rect 195686 453818 195728 454054
rect 195408 453734 195728 453818
rect 195408 453498 195450 453734
rect 195686 453498 195728 453734
rect 195408 453466 195728 453498
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 190288 414334 190608 414366
rect 190288 414098 190330 414334
rect 190566 414098 190608 414334
rect 190288 414014 190608 414098
rect 190288 413778 190330 414014
rect 190566 413778 190608 414014
rect 190288 413746 190608 413778
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 185168 374614 185488 374646
rect 185168 374378 185210 374614
rect 185446 374378 185488 374614
rect 185168 374294 185488 374378
rect 185168 374058 185210 374294
rect 185446 374058 185488 374294
rect 185168 374026 185488 374058
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 180048 334894 180368 334926
rect 180048 334658 180090 334894
rect 180326 334658 180368 334894
rect 180048 334574 180368 334658
rect 180048 334338 180090 334574
rect 180326 334338 180368 334574
rect 180048 334306 180368 334338
rect 174928 331174 175248 331206
rect 174928 330938 174970 331174
rect 175206 330938 175248 331174
rect 174928 330854 175248 330938
rect 174928 330618 174970 330854
rect 175206 330618 175248 330854
rect 174928 330586 175248 330618
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 169808 291454 170128 291486
rect 169808 291218 169850 291454
rect 170086 291218 170128 291454
rect 169808 291134 170128 291218
rect 169808 290898 169850 291134
rect 170086 290898 170128 291134
rect 169808 290866 170128 290898
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 164688 274054 165008 274086
rect 164688 273818 164730 274054
rect 164966 273818 165008 274054
rect 164688 273734 165008 273818
rect 164688 273498 164730 273734
rect 164966 273498 165008 273734
rect 164688 273466 165008 273498
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 133968 238054 134288 238086
rect 133968 237818 134010 238054
rect 134246 237818 134288 238054
rect 133968 237734 134288 237818
rect 133968 237498 134010 237734
rect 134246 237498 134288 237734
rect 133968 237466 134288 237498
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 113488 187174 113808 187206
rect 113488 186938 113530 187174
rect 113766 186938 113808 187174
rect 113488 186854 113808 186938
rect 113488 186618 113530 186854
rect 113766 186618 113808 186854
rect 113488 186586 113808 186618
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 99834 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 100454 173494
rect 99834 173174 100454 173258
rect 99834 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 100454 173174
rect 98128 162334 98448 162366
rect 98128 162098 98170 162334
rect 98406 162098 98448 162334
rect 98128 162014 98448 162098
rect 98128 161778 98170 162014
rect 98406 161778 98448 162014
rect 98128 161746 98448 161778
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 93008 122614 93328 122646
rect 93008 122378 93050 122614
rect 93286 122378 93328 122614
rect 93008 122294 93328 122378
rect 93008 122058 93050 122294
rect 93286 122058 93328 122294
rect 93008 122026 93328 122058
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 87888 82894 88208 82926
rect 87888 82658 87930 82894
rect 88166 82658 88208 82894
rect 87888 82574 88208 82658
rect 87888 82338 87930 82574
rect 88166 82338 88208 82574
rect 87888 82306 88208 82338
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 82768 43174 83088 43206
rect 82768 42938 82810 43174
rect 83046 42938 83088 43174
rect 82768 42854 83088 42938
rect 82768 42618 82810 42854
rect 83046 42618 83088 42854
rect 82768 42586 83088 42618
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 -1306 78134 2988
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 -2266 81854 10338
rect 84954 14614 85574 50058
rect 88674 54334 89294 89778
rect 96114 97774 96734 133218
rect 99834 137494 100454 172938
rect 103248 166054 103568 166086
rect 103248 165818 103290 166054
rect 103526 165818 103568 166054
rect 103248 165734 103568 165818
rect 103248 165498 103290 165734
rect 103526 165498 103568 165734
rect 103248 165466 103568 165498
rect 108368 147454 108688 147486
rect 108368 147218 108410 147454
rect 108646 147218 108688 147454
rect 108368 147134 108688 147218
rect 108368 146898 108410 147134
rect 108646 146898 108688 147134
rect 108368 146866 108688 146898
rect 109794 147454 110414 182898
rect 117234 154894 117854 190338
rect 118608 190894 118928 190926
rect 118608 190658 118650 190894
rect 118886 190658 118928 190894
rect 118608 190574 118928 190658
rect 118608 190338 118650 190574
rect 118886 190338 118928 190574
rect 118608 190306 118928 190338
rect 120954 158614 121574 194058
rect 123728 194614 124048 194646
rect 123728 194378 123770 194614
rect 124006 194378 124048 194614
rect 123728 194294 124048 194378
rect 123728 194058 123770 194294
rect 124006 194058 124048 194294
rect 123728 194026 124048 194058
rect 124674 162334 125294 197778
rect 128848 198334 129168 198366
rect 128848 198098 128890 198334
rect 129126 198098 129168 198334
rect 128848 198014 129168 198098
rect 128848 197778 128890 198014
rect 129126 197778 129168 198014
rect 128848 197746 129168 197778
rect 132114 169774 132734 205218
rect 135834 209494 136454 244938
rect 144208 223174 144528 223206
rect 144208 222938 144250 223174
rect 144486 222938 144528 223174
rect 144208 222854 144528 222938
rect 144208 222618 144250 222854
rect 144486 222618 144528 222854
rect 144208 222586 144528 222618
rect 139088 219454 139408 219486
rect 139088 219218 139130 219454
rect 139366 219218 139408 219454
rect 139088 219134 139408 219218
rect 139088 218898 139130 219134
rect 139366 218898 139408 219134
rect 139088 218866 139408 218898
rect 145794 219454 146414 254898
rect 149328 226894 149648 226926
rect 149328 226658 149370 226894
rect 149606 226658 149648 226894
rect 149328 226574 149648 226658
rect 149328 226338 149370 226574
rect 149606 226338 149648 226574
rect 149328 226306 149648 226338
rect 153234 226894 153854 262338
rect 154448 230614 154768 230646
rect 154448 230378 154490 230614
rect 154726 230378 154768 230614
rect 154448 230294 154768 230378
rect 154448 230058 154490 230294
rect 154726 230058 154768 230294
rect 154448 230026 154768 230058
rect 156954 230614 157574 266058
rect 159568 234334 159888 234366
rect 159568 234098 159610 234334
rect 159846 234098 159888 234334
rect 159568 234014 159888 234098
rect 159568 233778 159610 234014
rect 159846 233778 159888 234014
rect 159568 233746 159888 233778
rect 160674 234334 161294 269778
rect 168114 241774 168734 277218
rect 171834 281494 172454 316938
rect 181794 327454 182414 362898
rect 189234 370894 189854 406338
rect 192954 410614 193574 446058
rect 196674 450334 197294 485778
rect 204114 493774 204734 529218
rect 207834 533494 208454 568938
rect 217794 579454 218414 614898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221008 594334 221328 594366
rect 221008 594098 221050 594334
rect 221286 594098 221328 594334
rect 221008 594014 221328 594098
rect 221008 593778 221050 594014
rect 221286 593778 221328 594014
rect 221008 593746 221328 593778
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 215888 554614 216208 554646
rect 215888 554378 215930 554614
rect 216166 554378 216208 554614
rect 215888 554294 216208 554378
rect 215888 554058 215930 554294
rect 216166 554058 216208 554294
rect 215888 554026 216208 554058
rect 210768 550894 211088 550926
rect 210768 550658 210810 550894
rect 211046 550658 211088 550894
rect 210768 550574 211088 550658
rect 210768 550338 210810 550574
rect 211046 550338 211088 550574
rect 210768 550306 211088 550338
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 205648 511174 205968 511206
rect 205648 510938 205690 511174
rect 205926 510938 205968 511174
rect 205648 510854 205968 510938
rect 205648 510618 205690 510854
rect 205926 510618 205968 510854
rect 205648 510586 205968 510618
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 200528 471454 200848 471486
rect 200528 471218 200570 471454
rect 200806 471218 200848 471454
rect 200528 471134 200848 471218
rect 200528 470898 200570 471134
rect 200806 470898 200848 471134
rect 200528 470866 200848 470898
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 195408 418054 195728 418086
rect 195408 417818 195450 418054
rect 195686 417818 195728 418054
rect 195408 417734 195728 417818
rect 195408 417498 195450 417734
rect 195686 417498 195728 417734
rect 195408 417466 195728 417498
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 190288 378334 190608 378366
rect 190288 378098 190330 378334
rect 190566 378098 190608 378334
rect 190288 378014 190608 378098
rect 190288 377778 190330 378014
rect 190566 377778 190608 378014
rect 190288 377746 190608 377778
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 185168 338614 185488 338646
rect 185168 338378 185210 338614
rect 185446 338378 185488 338614
rect 185168 338294 185488 338378
rect 185168 338058 185210 338294
rect 185446 338058 185488 338294
rect 185168 338026 185488 338058
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 180048 298894 180368 298926
rect 180048 298658 180090 298894
rect 180326 298658 180368 298894
rect 180048 298574 180368 298658
rect 180048 298338 180090 298574
rect 180326 298338 180368 298574
rect 180048 298306 180368 298338
rect 174928 295174 175248 295206
rect 174928 294938 174970 295174
rect 175206 294938 175248 295174
rect 174928 294854 175248 294938
rect 174928 294618 174970 294854
rect 175206 294618 175248 294854
rect 174928 294586 175248 294618
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 169808 255454 170128 255486
rect 169808 255218 169850 255454
rect 170086 255218 170128 255454
rect 169808 255134 170128 255218
rect 169808 254898 169850 255134
rect 170086 254898 170128 255134
rect 169808 254866 170128 254898
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 164688 238054 165008 238086
rect 164688 237818 164730 238054
rect 164966 237818 165008 238054
rect 164688 237734 165008 237818
rect 164688 237498 164730 237734
rect 164966 237498 165008 237734
rect 164688 237466 165008 237498
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 133968 202054 134288 202086
rect 133968 201818 134010 202054
rect 134246 201818 134288 202054
rect 133968 201734 134288 201818
rect 133968 201498 134010 201734
rect 134246 201498 134288 201734
rect 133968 201466 134288 201498
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 113488 151174 113808 151206
rect 113488 150938 113530 151174
rect 113766 150938 113808 151174
rect 113488 150854 113808 150938
rect 113488 150618 113530 150854
rect 113766 150618 113808 150854
rect 113488 150586 113808 150618
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 99834 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 100454 137494
rect 99834 137174 100454 137258
rect 99834 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 100454 137174
rect 98128 126334 98448 126366
rect 98128 126098 98170 126334
rect 98406 126098 98448 126334
rect 98128 126014 98448 126098
rect 98128 125778 98170 126014
rect 98406 125778 98448 126014
rect 98128 125746 98448 125778
rect 96114 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 96734 97774
rect 96114 97454 96734 97538
rect 96114 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 96734 97454
rect 93008 86614 93328 86646
rect 93008 86378 93050 86614
rect 93286 86378 93328 86614
rect 93008 86294 93328 86378
rect 93008 86058 93050 86294
rect 93286 86058 93328 86294
rect 93008 86026 93328 86058
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 87888 46894 88208 46926
rect 87888 46658 87930 46894
rect 88166 46658 88208 46894
rect 87888 46574 88208 46658
rect 87888 46338 87930 46574
rect 88166 46338 88208 46574
rect 87888 46306 88208 46338
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 82768 7174 83088 7206
rect 82768 6938 82810 7174
rect 83046 6938 83088 7174
rect 82768 6854 83088 6938
rect 82768 6618 82810 6854
rect 83046 6618 83088 6854
rect 82768 6586 83088 6618
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 -3226 85574 14058
rect 88674 18334 89294 53778
rect 96114 61774 96734 97218
rect 99834 101494 100454 136938
rect 103248 130054 103568 130086
rect 103248 129818 103290 130054
rect 103526 129818 103568 130054
rect 103248 129734 103568 129818
rect 103248 129498 103290 129734
rect 103526 129498 103568 129734
rect 103248 129466 103568 129498
rect 108368 111454 108688 111486
rect 108368 111218 108410 111454
rect 108646 111218 108688 111454
rect 108368 111134 108688 111218
rect 108368 110898 108410 111134
rect 108646 110898 108688 111134
rect 108368 110866 108688 110898
rect 109794 111454 110414 146898
rect 117234 118894 117854 154338
rect 118608 154894 118928 154926
rect 118608 154658 118650 154894
rect 118886 154658 118928 154894
rect 118608 154574 118928 154658
rect 118608 154338 118650 154574
rect 118886 154338 118928 154574
rect 118608 154306 118928 154338
rect 120954 122614 121574 158058
rect 123728 158614 124048 158646
rect 123728 158378 123770 158614
rect 124006 158378 124048 158614
rect 123728 158294 124048 158378
rect 123728 158058 123770 158294
rect 124006 158058 124048 158294
rect 123728 158026 124048 158058
rect 124674 126334 125294 161778
rect 128848 162334 129168 162366
rect 128848 162098 128890 162334
rect 129126 162098 129168 162334
rect 128848 162014 129168 162098
rect 128848 161778 128890 162014
rect 129126 161778 129168 162014
rect 128848 161746 129168 161778
rect 132114 133774 132734 169218
rect 135834 173494 136454 208938
rect 144208 187174 144528 187206
rect 144208 186938 144250 187174
rect 144486 186938 144528 187174
rect 144208 186854 144528 186938
rect 144208 186618 144250 186854
rect 144486 186618 144528 186854
rect 144208 186586 144528 186618
rect 139088 183454 139408 183486
rect 139088 183218 139130 183454
rect 139366 183218 139408 183454
rect 139088 183134 139408 183218
rect 139088 182898 139130 183134
rect 139366 182898 139408 183134
rect 139088 182866 139408 182898
rect 145794 183454 146414 218898
rect 149328 190894 149648 190926
rect 149328 190658 149370 190894
rect 149606 190658 149648 190894
rect 149328 190574 149648 190658
rect 149328 190338 149370 190574
rect 149606 190338 149648 190574
rect 149328 190306 149648 190338
rect 153234 190894 153854 226338
rect 154448 194614 154768 194646
rect 154448 194378 154490 194614
rect 154726 194378 154768 194614
rect 154448 194294 154768 194378
rect 154448 194058 154490 194294
rect 154726 194058 154768 194294
rect 154448 194026 154768 194058
rect 156954 194614 157574 230058
rect 159568 198334 159888 198366
rect 159568 198098 159610 198334
rect 159846 198098 159888 198334
rect 159568 198014 159888 198098
rect 159568 197778 159610 198014
rect 159846 197778 159888 198014
rect 159568 197746 159888 197778
rect 160674 198334 161294 233778
rect 168114 205774 168734 241218
rect 171834 245494 172454 280938
rect 181794 291454 182414 326898
rect 189234 334894 189854 370338
rect 192954 374614 193574 410058
rect 196674 414334 197294 449778
rect 204114 457774 204734 493218
rect 207834 497494 208454 532938
rect 217794 543454 218414 578898
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221008 558334 221328 558366
rect 221008 558098 221050 558334
rect 221286 558098 221328 558334
rect 221008 558014 221328 558098
rect 221008 557778 221050 558014
rect 221286 557778 221328 558014
rect 221008 557746 221328 557778
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 215888 518614 216208 518646
rect 215888 518378 215930 518614
rect 216166 518378 216208 518614
rect 215888 518294 216208 518378
rect 215888 518058 215930 518294
rect 216166 518058 216208 518294
rect 215888 518026 216208 518058
rect 210768 514894 211088 514926
rect 210768 514658 210810 514894
rect 211046 514658 211088 514894
rect 210768 514574 211088 514658
rect 210768 514338 210810 514574
rect 211046 514338 211088 514574
rect 210768 514306 211088 514338
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 205648 475174 205968 475206
rect 205648 474938 205690 475174
rect 205926 474938 205968 475174
rect 205648 474854 205968 474938
rect 205648 474618 205690 474854
rect 205926 474618 205968 474854
rect 205648 474586 205968 474618
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 200528 435454 200848 435486
rect 200528 435218 200570 435454
rect 200806 435218 200848 435454
rect 200528 435134 200848 435218
rect 200528 434898 200570 435134
rect 200806 434898 200848 435134
rect 200528 434866 200848 434898
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 195408 382054 195728 382086
rect 195408 381818 195450 382054
rect 195686 381818 195728 382054
rect 195408 381734 195728 381818
rect 195408 381498 195450 381734
rect 195686 381498 195728 381734
rect 195408 381466 195728 381498
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 190288 342334 190608 342366
rect 190288 342098 190330 342334
rect 190566 342098 190608 342334
rect 190288 342014 190608 342098
rect 190288 341778 190330 342014
rect 190566 341778 190608 342014
rect 190288 341746 190608 341778
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 185168 302614 185488 302646
rect 185168 302378 185210 302614
rect 185446 302378 185488 302614
rect 185168 302294 185488 302378
rect 185168 302058 185210 302294
rect 185446 302058 185488 302294
rect 185168 302026 185488 302058
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 180048 262894 180368 262926
rect 180048 262658 180090 262894
rect 180326 262658 180368 262894
rect 180048 262574 180368 262658
rect 180048 262338 180090 262574
rect 180326 262338 180368 262574
rect 180048 262306 180368 262338
rect 174928 259174 175248 259206
rect 174928 258938 174970 259174
rect 175206 258938 175248 259174
rect 174928 258854 175248 258938
rect 174928 258618 174970 258854
rect 175206 258618 175248 258854
rect 174928 258586 175248 258618
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 169808 219454 170128 219486
rect 169808 219218 169850 219454
rect 170086 219218 170128 219454
rect 169808 219134 170128 219218
rect 169808 218898 169850 219134
rect 170086 218898 170128 219134
rect 169808 218866 170128 218898
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 164688 202054 165008 202086
rect 164688 201818 164730 202054
rect 164966 201818 165008 202054
rect 164688 201734 165008 201818
rect 164688 201498 164730 201734
rect 164966 201498 165008 201734
rect 164688 201466 165008 201498
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 133968 166054 134288 166086
rect 133968 165818 134010 166054
rect 134246 165818 134288 166054
rect 133968 165734 134288 165818
rect 133968 165498 134010 165734
rect 134246 165498 134288 165734
rect 133968 165466 134288 165498
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 113488 115174 113808 115206
rect 113488 114938 113530 115174
rect 113766 114938 113808 115174
rect 113488 114854 113808 114938
rect 113488 114618 113530 114854
rect 113766 114618 113808 114854
rect 113488 114586 113808 114618
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 99834 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 100454 101494
rect 99834 101174 100454 101258
rect 99834 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 100454 101174
rect 98128 90334 98448 90366
rect 98128 90098 98170 90334
rect 98406 90098 98448 90334
rect 98128 90014 98448 90098
rect 98128 89778 98170 90014
rect 98406 89778 98448 90014
rect 98128 89746 98448 89778
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 93008 50614 93328 50646
rect 93008 50378 93050 50614
rect 93286 50378 93328 50614
rect 93008 50294 93328 50378
rect 93008 50058 93050 50294
rect 93286 50058 93328 50294
rect 93008 50026 93328 50058
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 87888 10894 88208 10926
rect 87888 10658 87930 10894
rect 88166 10658 88208 10894
rect 87888 10574 88208 10658
rect 87888 10338 87930 10574
rect 88166 10338 88208 10574
rect 87888 10306 88208 10338
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 -4186 89294 17778
rect 96114 25774 96734 61218
rect 99834 65494 100454 100938
rect 103248 94054 103568 94086
rect 103248 93818 103290 94054
rect 103526 93818 103568 94054
rect 103248 93734 103568 93818
rect 103248 93498 103290 93734
rect 103526 93498 103568 93734
rect 103248 93466 103568 93498
rect 108368 75454 108688 75486
rect 108368 75218 108410 75454
rect 108646 75218 108688 75454
rect 108368 75134 108688 75218
rect 108368 74898 108410 75134
rect 108646 74898 108688 75134
rect 108368 74866 108688 74898
rect 109794 75454 110414 110898
rect 117234 82894 117854 118338
rect 118608 118894 118928 118926
rect 118608 118658 118650 118894
rect 118886 118658 118928 118894
rect 118608 118574 118928 118658
rect 118608 118338 118650 118574
rect 118886 118338 118928 118574
rect 118608 118306 118928 118338
rect 120954 86614 121574 122058
rect 123728 122614 124048 122646
rect 123728 122378 123770 122614
rect 124006 122378 124048 122614
rect 123728 122294 124048 122378
rect 123728 122058 123770 122294
rect 124006 122058 124048 122294
rect 123728 122026 124048 122058
rect 124674 90334 125294 125778
rect 128848 126334 129168 126366
rect 128848 126098 128890 126334
rect 129126 126098 129168 126334
rect 128848 126014 129168 126098
rect 128848 125778 128890 126014
rect 129126 125778 129168 126014
rect 128848 125746 129168 125778
rect 132114 97774 132734 133218
rect 135834 137494 136454 172938
rect 144208 151174 144528 151206
rect 144208 150938 144250 151174
rect 144486 150938 144528 151174
rect 144208 150854 144528 150938
rect 144208 150618 144250 150854
rect 144486 150618 144528 150854
rect 144208 150586 144528 150618
rect 139088 147454 139408 147486
rect 139088 147218 139130 147454
rect 139366 147218 139408 147454
rect 139088 147134 139408 147218
rect 139088 146898 139130 147134
rect 139366 146898 139408 147134
rect 139088 146866 139408 146898
rect 145794 147454 146414 182898
rect 149328 154894 149648 154926
rect 149328 154658 149370 154894
rect 149606 154658 149648 154894
rect 149328 154574 149648 154658
rect 149328 154338 149370 154574
rect 149606 154338 149648 154574
rect 149328 154306 149648 154338
rect 153234 154894 153854 190338
rect 154448 158614 154768 158646
rect 154448 158378 154490 158614
rect 154726 158378 154768 158614
rect 154448 158294 154768 158378
rect 154448 158058 154490 158294
rect 154726 158058 154768 158294
rect 154448 158026 154768 158058
rect 156954 158614 157574 194058
rect 159568 162334 159888 162366
rect 159568 162098 159610 162334
rect 159846 162098 159888 162334
rect 159568 162014 159888 162098
rect 159568 161778 159610 162014
rect 159846 161778 159888 162014
rect 159568 161746 159888 161778
rect 160674 162334 161294 197778
rect 168114 169774 168734 205218
rect 171834 209494 172454 244938
rect 181794 255454 182414 290898
rect 189234 298894 189854 334338
rect 192954 338614 193574 374058
rect 196674 378334 197294 413778
rect 204114 421774 204734 457218
rect 207834 461494 208454 496938
rect 217794 507454 218414 542898
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221008 522334 221328 522366
rect 221008 522098 221050 522334
rect 221286 522098 221328 522334
rect 221008 522014 221328 522098
rect 221008 521778 221050 522014
rect 221286 521778 221328 522014
rect 221008 521746 221328 521778
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 215888 482614 216208 482646
rect 215888 482378 215930 482614
rect 216166 482378 216208 482614
rect 215888 482294 216208 482378
rect 215888 482058 215930 482294
rect 216166 482058 216208 482294
rect 215888 482026 216208 482058
rect 210768 478894 211088 478926
rect 210768 478658 210810 478894
rect 211046 478658 211088 478894
rect 210768 478574 211088 478658
rect 210768 478338 210810 478574
rect 211046 478338 211088 478574
rect 210768 478306 211088 478338
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 205648 439174 205968 439206
rect 205648 438938 205690 439174
rect 205926 438938 205968 439174
rect 205648 438854 205968 438938
rect 205648 438618 205690 438854
rect 205926 438618 205968 438854
rect 205648 438586 205968 438618
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 200528 399454 200848 399486
rect 200528 399218 200570 399454
rect 200806 399218 200848 399454
rect 200528 399134 200848 399218
rect 200528 398898 200570 399134
rect 200806 398898 200848 399134
rect 200528 398866 200848 398898
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 195408 346054 195728 346086
rect 195408 345818 195450 346054
rect 195686 345818 195728 346054
rect 195408 345734 195728 345818
rect 195408 345498 195450 345734
rect 195686 345498 195728 345734
rect 195408 345466 195728 345498
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 190288 306334 190608 306366
rect 190288 306098 190330 306334
rect 190566 306098 190608 306334
rect 190288 306014 190608 306098
rect 190288 305778 190330 306014
rect 190566 305778 190608 306014
rect 190288 305746 190608 305778
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 185168 266614 185488 266646
rect 185168 266378 185210 266614
rect 185446 266378 185488 266614
rect 185168 266294 185488 266378
rect 185168 266058 185210 266294
rect 185446 266058 185488 266294
rect 185168 266026 185488 266058
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 180048 226894 180368 226926
rect 180048 226658 180090 226894
rect 180326 226658 180368 226894
rect 180048 226574 180368 226658
rect 180048 226338 180090 226574
rect 180326 226338 180368 226574
rect 180048 226306 180368 226338
rect 174928 223174 175248 223206
rect 174928 222938 174970 223174
rect 175206 222938 175248 223174
rect 174928 222854 175248 222938
rect 174928 222618 174970 222854
rect 175206 222618 175248 222854
rect 174928 222586 175248 222618
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 169808 183454 170128 183486
rect 169808 183218 169850 183454
rect 170086 183218 170128 183454
rect 169808 183134 170128 183218
rect 169808 182898 169850 183134
rect 170086 182898 170128 183134
rect 169808 182866 170128 182898
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 164688 166054 165008 166086
rect 164688 165818 164730 166054
rect 164966 165818 165008 166054
rect 164688 165734 165008 165818
rect 164688 165498 164730 165734
rect 164966 165498 165008 165734
rect 164688 165466 165008 165498
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 133968 130054 134288 130086
rect 133968 129818 134010 130054
rect 134246 129818 134288 130054
rect 133968 129734 134288 129818
rect 133968 129498 134010 129734
rect 134246 129498 134288 129734
rect 133968 129466 134288 129498
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 113488 79174 113808 79206
rect 113488 78938 113530 79174
rect 113766 78938 113808 79174
rect 113488 78854 113808 78938
rect 113488 78618 113530 78854
rect 113766 78618 113808 78854
rect 113488 78586 113808 78618
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 98128 54334 98448 54366
rect 98128 54098 98170 54334
rect 98406 54098 98448 54334
rect 98128 54014 98448 54098
rect 98128 53778 98170 54014
rect 98406 53778 98448 54014
rect 98128 53746 98448 53778
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 93008 14614 93328 14646
rect 93008 14378 93050 14614
rect 93286 14378 93328 14614
rect 93008 14294 93328 14378
rect 93008 14058 93050 14294
rect 93286 14058 93328 14294
rect 93008 14026 93328 14058
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 -5146 93014 2988
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 -6106 96734 25218
rect 99834 29494 100454 64938
rect 103248 58054 103568 58086
rect 103248 57818 103290 58054
rect 103526 57818 103568 58054
rect 103248 57734 103568 57818
rect 103248 57498 103290 57734
rect 103526 57498 103568 57734
rect 103248 57466 103568 57498
rect 108368 39454 108688 39486
rect 108368 39218 108410 39454
rect 108646 39218 108688 39454
rect 108368 39134 108688 39218
rect 108368 38898 108410 39134
rect 108646 38898 108688 39134
rect 108368 38866 108688 38898
rect 109794 39454 110414 74898
rect 117234 46894 117854 82338
rect 118608 82894 118928 82926
rect 118608 82658 118650 82894
rect 118886 82658 118928 82894
rect 118608 82574 118928 82658
rect 118608 82338 118650 82574
rect 118886 82338 118928 82574
rect 118608 82306 118928 82338
rect 120954 50614 121574 86058
rect 123728 86614 124048 86646
rect 123728 86378 123770 86614
rect 124006 86378 124048 86614
rect 123728 86294 124048 86378
rect 123728 86058 123770 86294
rect 124006 86058 124048 86294
rect 123728 86026 124048 86058
rect 124674 54334 125294 89778
rect 128848 90334 129168 90366
rect 128848 90098 128890 90334
rect 129126 90098 129168 90334
rect 128848 90014 129168 90098
rect 128848 89778 128890 90014
rect 129126 89778 129168 90014
rect 128848 89746 129168 89778
rect 132114 61774 132734 97218
rect 135834 101494 136454 136938
rect 144208 115174 144528 115206
rect 144208 114938 144250 115174
rect 144486 114938 144528 115174
rect 144208 114854 144528 114938
rect 144208 114618 144250 114854
rect 144486 114618 144528 114854
rect 144208 114586 144528 114618
rect 139088 111454 139408 111486
rect 139088 111218 139130 111454
rect 139366 111218 139408 111454
rect 139088 111134 139408 111218
rect 139088 110898 139130 111134
rect 139366 110898 139408 111134
rect 139088 110866 139408 110898
rect 145794 111454 146414 146898
rect 149328 118894 149648 118926
rect 149328 118658 149370 118894
rect 149606 118658 149648 118894
rect 149328 118574 149648 118658
rect 149328 118338 149370 118574
rect 149606 118338 149648 118574
rect 149328 118306 149648 118338
rect 153234 118894 153854 154338
rect 154448 122614 154768 122646
rect 154448 122378 154490 122614
rect 154726 122378 154768 122614
rect 154448 122294 154768 122378
rect 154448 122058 154490 122294
rect 154726 122058 154768 122294
rect 154448 122026 154768 122058
rect 156954 122614 157574 158058
rect 159568 126334 159888 126366
rect 159568 126098 159610 126334
rect 159846 126098 159888 126334
rect 159568 126014 159888 126098
rect 159568 125778 159610 126014
rect 159846 125778 159888 126014
rect 159568 125746 159888 125778
rect 160674 126334 161294 161778
rect 168114 133774 168734 169218
rect 171834 173494 172454 208938
rect 181794 219454 182414 254898
rect 189234 262894 189854 298338
rect 192954 302614 193574 338058
rect 196674 342334 197294 377778
rect 204114 385774 204734 421218
rect 207834 425494 208454 460938
rect 217794 471454 218414 506898
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221008 486334 221328 486366
rect 221008 486098 221050 486334
rect 221286 486098 221328 486334
rect 221008 486014 221328 486098
rect 221008 485778 221050 486014
rect 221286 485778 221328 486014
rect 221008 485746 221328 485778
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 215888 446614 216208 446646
rect 215888 446378 215930 446614
rect 216166 446378 216208 446614
rect 215888 446294 216208 446378
rect 215888 446058 215930 446294
rect 216166 446058 216208 446294
rect 215888 446026 216208 446058
rect 210768 442894 211088 442926
rect 210768 442658 210810 442894
rect 211046 442658 211088 442894
rect 210768 442574 211088 442658
rect 210768 442338 210810 442574
rect 211046 442338 211088 442574
rect 210768 442306 211088 442338
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 205648 403174 205968 403206
rect 205648 402938 205690 403174
rect 205926 402938 205968 403174
rect 205648 402854 205968 402938
rect 205648 402618 205690 402854
rect 205926 402618 205968 402854
rect 205648 402586 205968 402618
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 200528 363454 200848 363486
rect 200528 363218 200570 363454
rect 200806 363218 200848 363454
rect 200528 363134 200848 363218
rect 200528 362898 200570 363134
rect 200806 362898 200848 363134
rect 200528 362866 200848 362898
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 195408 310054 195728 310086
rect 195408 309818 195450 310054
rect 195686 309818 195728 310054
rect 195408 309734 195728 309818
rect 195408 309498 195450 309734
rect 195686 309498 195728 309734
rect 195408 309466 195728 309498
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 190288 270334 190608 270366
rect 190288 270098 190330 270334
rect 190566 270098 190608 270334
rect 190288 270014 190608 270098
rect 190288 269778 190330 270014
rect 190566 269778 190608 270014
rect 190288 269746 190608 269778
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 185168 230614 185488 230646
rect 185168 230378 185210 230614
rect 185446 230378 185488 230614
rect 185168 230294 185488 230378
rect 185168 230058 185210 230294
rect 185446 230058 185488 230294
rect 185168 230026 185488 230058
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 180048 190894 180368 190926
rect 180048 190658 180090 190894
rect 180326 190658 180368 190894
rect 180048 190574 180368 190658
rect 180048 190338 180090 190574
rect 180326 190338 180368 190574
rect 180048 190306 180368 190338
rect 174928 187174 175248 187206
rect 174928 186938 174970 187174
rect 175206 186938 175248 187174
rect 174928 186854 175248 186938
rect 174928 186618 174970 186854
rect 175206 186618 175248 186854
rect 174928 186586 175248 186618
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 169808 147454 170128 147486
rect 169808 147218 169850 147454
rect 170086 147218 170128 147454
rect 169808 147134 170128 147218
rect 169808 146898 169850 147134
rect 170086 146898 170128 147134
rect 169808 146866 170128 146898
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 164688 130054 165008 130086
rect 164688 129818 164730 130054
rect 164966 129818 165008 130054
rect 164688 129734 165008 129818
rect 164688 129498 164730 129734
rect 164966 129498 165008 129734
rect 164688 129466 165008 129498
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 133968 94054 134288 94086
rect 133968 93818 134010 94054
rect 134246 93818 134288 94054
rect 133968 93734 134288 93818
rect 133968 93498 134010 93734
rect 134246 93498 134288 93734
rect 133968 93466 134288 93498
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 113488 43174 113808 43206
rect 113488 42938 113530 43174
rect 113766 42938 113808 43174
rect 113488 42854 113808 42938
rect 113488 42618 113530 42854
rect 113766 42618 113808 42854
rect 113488 42586 113808 42618
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 98128 18334 98448 18366
rect 98128 18098 98170 18334
rect 98406 18098 98448 18334
rect 98128 18014 98448 18098
rect 98128 17778 98170 18014
rect 98406 17778 98448 18014
rect 98128 17746 98448 17778
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 -7066 100454 28938
rect 103248 22054 103568 22086
rect 103248 21818 103290 22054
rect 103526 21818 103568 22054
rect 103248 21734 103568 21818
rect 103248 21498 103290 21734
rect 103526 21498 103568 21734
rect 103248 21466 103568 21498
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 3454 110414 38898
rect 117234 10894 117854 46338
rect 118608 46894 118928 46926
rect 118608 46658 118650 46894
rect 118886 46658 118928 46894
rect 118608 46574 118928 46658
rect 118608 46338 118650 46574
rect 118886 46338 118928 46574
rect 118608 46306 118928 46338
rect 120954 14614 121574 50058
rect 123728 50614 124048 50646
rect 123728 50378 123770 50614
rect 124006 50378 124048 50614
rect 123728 50294 124048 50378
rect 123728 50058 123770 50294
rect 124006 50058 124048 50294
rect 123728 50026 124048 50058
rect 124674 18334 125294 53778
rect 128848 54334 129168 54366
rect 128848 54098 128890 54334
rect 129126 54098 129168 54334
rect 128848 54014 129168 54098
rect 128848 53778 128890 54014
rect 129126 53778 129168 54014
rect 128848 53746 129168 53778
rect 132114 25774 132734 61218
rect 135834 65494 136454 100938
rect 144208 79174 144528 79206
rect 144208 78938 144250 79174
rect 144486 78938 144528 79174
rect 144208 78854 144528 78938
rect 144208 78618 144250 78854
rect 144486 78618 144528 78854
rect 144208 78586 144528 78618
rect 139088 75454 139408 75486
rect 139088 75218 139130 75454
rect 139366 75218 139408 75454
rect 139088 75134 139408 75218
rect 139088 74898 139130 75134
rect 139366 74898 139408 75134
rect 139088 74866 139408 74898
rect 145794 75454 146414 110898
rect 149328 82894 149648 82926
rect 149328 82658 149370 82894
rect 149606 82658 149648 82894
rect 149328 82574 149648 82658
rect 149328 82338 149370 82574
rect 149606 82338 149648 82574
rect 149328 82306 149648 82338
rect 153234 82894 153854 118338
rect 154448 86614 154768 86646
rect 154448 86378 154490 86614
rect 154726 86378 154768 86614
rect 154448 86294 154768 86378
rect 154448 86058 154490 86294
rect 154726 86058 154768 86294
rect 154448 86026 154768 86058
rect 156954 86614 157574 122058
rect 159568 90334 159888 90366
rect 159568 90098 159610 90334
rect 159846 90098 159888 90334
rect 159568 90014 159888 90098
rect 159568 89778 159610 90014
rect 159846 89778 159888 90014
rect 159568 89746 159888 89778
rect 160674 90334 161294 125778
rect 168114 97774 168734 133218
rect 171834 137494 172454 172938
rect 181794 183454 182414 218898
rect 189234 226894 189854 262338
rect 192954 266614 193574 302058
rect 196674 306334 197294 341778
rect 204114 349774 204734 385218
rect 207834 389494 208454 424938
rect 217794 435454 218414 470898
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221008 450334 221328 450366
rect 221008 450098 221050 450334
rect 221286 450098 221328 450334
rect 221008 450014 221328 450098
rect 221008 449778 221050 450014
rect 221286 449778 221328 450014
rect 221008 449746 221328 449778
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 215888 410614 216208 410646
rect 215888 410378 215930 410614
rect 216166 410378 216208 410614
rect 215888 410294 216208 410378
rect 215888 410058 215930 410294
rect 216166 410058 216208 410294
rect 215888 410026 216208 410058
rect 210768 406894 211088 406926
rect 210768 406658 210810 406894
rect 211046 406658 211088 406894
rect 210768 406574 211088 406658
rect 210768 406338 210810 406574
rect 211046 406338 211088 406574
rect 210768 406306 211088 406338
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 205648 367174 205968 367206
rect 205648 366938 205690 367174
rect 205926 366938 205968 367174
rect 205648 366854 205968 366938
rect 205648 366618 205690 366854
rect 205926 366618 205968 366854
rect 205648 366586 205968 366618
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 200528 327454 200848 327486
rect 200528 327218 200570 327454
rect 200806 327218 200848 327454
rect 200528 327134 200848 327218
rect 200528 326898 200570 327134
rect 200806 326898 200848 327134
rect 200528 326866 200848 326898
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 195408 274054 195728 274086
rect 195408 273818 195450 274054
rect 195686 273818 195728 274054
rect 195408 273734 195728 273818
rect 195408 273498 195450 273734
rect 195686 273498 195728 273734
rect 195408 273466 195728 273498
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 190288 234334 190608 234366
rect 190288 234098 190330 234334
rect 190566 234098 190608 234334
rect 190288 234014 190608 234098
rect 190288 233778 190330 234014
rect 190566 233778 190608 234014
rect 190288 233746 190608 233778
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 185168 194614 185488 194646
rect 185168 194378 185210 194614
rect 185446 194378 185488 194614
rect 185168 194294 185488 194378
rect 185168 194058 185210 194294
rect 185446 194058 185488 194294
rect 185168 194026 185488 194058
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 180048 154894 180368 154926
rect 180048 154658 180090 154894
rect 180326 154658 180368 154894
rect 180048 154574 180368 154658
rect 180048 154338 180090 154574
rect 180326 154338 180368 154574
rect 180048 154306 180368 154338
rect 174928 151174 175248 151206
rect 174928 150938 174970 151174
rect 175206 150938 175248 151174
rect 174928 150854 175248 150938
rect 174928 150618 174970 150854
rect 175206 150618 175248 150854
rect 174928 150586 175248 150618
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 169808 111454 170128 111486
rect 169808 111218 169850 111454
rect 170086 111218 170128 111454
rect 169808 111134 170128 111218
rect 169808 110898 169850 111134
rect 170086 110898 170128 111134
rect 169808 110866 170128 110898
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 164688 94054 165008 94086
rect 164688 93818 164730 94054
rect 164966 93818 165008 94054
rect 164688 93734 165008 93818
rect 164688 93498 164730 93734
rect 164966 93498 165008 93734
rect 164688 93466 165008 93498
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 133968 58054 134288 58086
rect 133968 57818 134010 58054
rect 134246 57818 134288 58054
rect 133968 57734 134288 57818
rect 133968 57498 134010 57734
rect 134246 57498 134288 57734
rect 133968 57466 134288 57498
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 113488 7174 113808 7206
rect 113488 6938 113530 7174
rect 113766 6938 113808 7174
rect 113488 6854 113808 6938
rect 113488 6618 113530 6854
rect 113766 6618 113808 6854
rect 113488 6586 113808 6618
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 -1306 114134 2988
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 -2266 117854 10338
rect 118608 10894 118928 10926
rect 118608 10658 118650 10894
rect 118886 10658 118928 10894
rect 118608 10574 118928 10658
rect 118608 10338 118650 10574
rect 118886 10338 118928 10574
rect 118608 10306 118928 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 -3226 121574 14058
rect 123728 14614 124048 14646
rect 123728 14378 123770 14614
rect 124006 14378 124048 14614
rect 123728 14294 124048 14378
rect 123728 14058 123770 14294
rect 124006 14058 124048 14294
rect 123728 14026 124048 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 -4186 125294 17778
rect 128848 18334 129168 18366
rect 128848 18098 128890 18334
rect 129126 18098 129168 18334
rect 128848 18014 129168 18098
rect 128848 17778 128890 18014
rect 129126 17778 129168 18014
rect 128848 17746 129168 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 -5146 129014 2988
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 -6106 132734 25218
rect 135834 29494 136454 64938
rect 144208 43174 144528 43206
rect 144208 42938 144250 43174
rect 144486 42938 144528 43174
rect 144208 42854 144528 42938
rect 144208 42618 144250 42854
rect 144486 42618 144528 42854
rect 144208 42586 144528 42618
rect 139088 39454 139408 39486
rect 139088 39218 139130 39454
rect 139366 39218 139408 39454
rect 139088 39134 139408 39218
rect 139088 38898 139130 39134
rect 139366 38898 139408 39134
rect 139088 38866 139408 38898
rect 145794 39454 146414 74898
rect 149328 46894 149648 46926
rect 149328 46658 149370 46894
rect 149606 46658 149648 46894
rect 149328 46574 149648 46658
rect 149328 46338 149370 46574
rect 149606 46338 149648 46574
rect 149328 46306 149648 46338
rect 153234 46894 153854 82338
rect 154448 50614 154768 50646
rect 154448 50378 154490 50614
rect 154726 50378 154768 50614
rect 154448 50294 154768 50378
rect 154448 50058 154490 50294
rect 154726 50058 154768 50294
rect 154448 50026 154768 50058
rect 156954 50614 157574 86058
rect 159568 54334 159888 54366
rect 159568 54098 159610 54334
rect 159846 54098 159888 54334
rect 159568 54014 159888 54098
rect 159568 53778 159610 54014
rect 159846 53778 159888 54014
rect 159568 53746 159888 53778
rect 160674 54334 161294 89778
rect 168114 61774 168734 97218
rect 171834 101494 172454 136938
rect 181794 147454 182414 182898
rect 189234 190894 189854 226338
rect 192954 230614 193574 266058
rect 196674 270334 197294 305778
rect 204114 313774 204734 349218
rect 207834 353494 208454 388938
rect 217794 399454 218414 434898
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221008 414334 221328 414366
rect 221008 414098 221050 414334
rect 221286 414098 221328 414334
rect 221008 414014 221328 414098
rect 221008 413778 221050 414014
rect 221286 413778 221328 414014
rect 221008 413746 221328 413778
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 215888 374614 216208 374646
rect 215888 374378 215930 374614
rect 216166 374378 216208 374614
rect 215888 374294 216208 374378
rect 215888 374058 215930 374294
rect 216166 374058 216208 374294
rect 215888 374026 216208 374058
rect 210768 370894 211088 370926
rect 210768 370658 210810 370894
rect 211046 370658 211088 370894
rect 210768 370574 211088 370658
rect 210768 370338 210810 370574
rect 211046 370338 211088 370574
rect 210768 370306 211088 370338
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 205648 331174 205968 331206
rect 205648 330938 205690 331174
rect 205926 330938 205968 331174
rect 205648 330854 205968 330938
rect 205648 330618 205690 330854
rect 205926 330618 205968 330854
rect 205648 330586 205968 330618
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 200528 291454 200848 291486
rect 200528 291218 200570 291454
rect 200806 291218 200848 291454
rect 200528 291134 200848 291218
rect 200528 290898 200570 291134
rect 200806 290898 200848 291134
rect 200528 290866 200848 290898
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 195408 238054 195728 238086
rect 195408 237818 195450 238054
rect 195686 237818 195728 238054
rect 195408 237734 195728 237818
rect 195408 237498 195450 237734
rect 195686 237498 195728 237734
rect 195408 237466 195728 237498
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 190288 198334 190608 198366
rect 190288 198098 190330 198334
rect 190566 198098 190608 198334
rect 190288 198014 190608 198098
rect 190288 197778 190330 198014
rect 190566 197778 190608 198014
rect 190288 197746 190608 197778
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 185168 158614 185488 158646
rect 185168 158378 185210 158614
rect 185446 158378 185488 158614
rect 185168 158294 185488 158378
rect 185168 158058 185210 158294
rect 185446 158058 185488 158294
rect 185168 158026 185488 158058
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 180048 118894 180368 118926
rect 180048 118658 180090 118894
rect 180326 118658 180368 118894
rect 180048 118574 180368 118658
rect 180048 118338 180090 118574
rect 180326 118338 180368 118574
rect 180048 118306 180368 118338
rect 174928 115174 175248 115206
rect 174928 114938 174970 115174
rect 175206 114938 175248 115174
rect 174928 114854 175248 114938
rect 174928 114618 174970 114854
rect 175206 114618 175248 114854
rect 174928 114586 175248 114618
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 169808 75454 170128 75486
rect 169808 75218 169850 75454
rect 170086 75218 170128 75454
rect 169808 75134 170128 75218
rect 169808 74898 169850 75134
rect 170086 74898 170128 75134
rect 169808 74866 170128 74898
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 164688 58054 165008 58086
rect 164688 57818 164730 58054
rect 164966 57818 165008 58054
rect 164688 57734 165008 57818
rect 164688 57498 164730 57734
rect 164966 57498 165008 57734
rect 164688 57466 165008 57498
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 133968 22054 134288 22086
rect 133968 21818 134010 22054
rect 134246 21818 134288 22054
rect 133968 21734 134288 21818
rect 133968 21498 134010 21734
rect 134246 21498 134288 21734
rect 133968 21466 134288 21498
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 -7066 136454 28938
rect 144208 7174 144528 7206
rect 144208 6938 144250 7174
rect 144486 6938 144528 7174
rect 144208 6854 144528 6938
rect 144208 6618 144250 6854
rect 144486 6618 144528 6854
rect 144208 6586 144528 6618
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 3454 146414 38898
rect 149328 10894 149648 10926
rect 149328 10658 149370 10894
rect 149606 10658 149648 10894
rect 149328 10574 149648 10658
rect 149328 10338 149370 10574
rect 149606 10338 149648 10574
rect 149328 10306 149648 10338
rect 153234 10894 153854 46338
rect 154448 14614 154768 14646
rect 154448 14378 154490 14614
rect 154726 14378 154768 14614
rect 154448 14294 154768 14378
rect 154448 14058 154490 14294
rect 154726 14058 154768 14294
rect 154448 14026 154768 14058
rect 156954 14614 157574 50058
rect 159568 18334 159888 18366
rect 159568 18098 159610 18334
rect 159846 18098 159888 18334
rect 159568 18014 159888 18098
rect 159568 17778 159610 18014
rect 159846 17778 159888 18014
rect 159568 17746 159888 17778
rect 160674 18334 161294 53778
rect 168114 25774 168734 61218
rect 171834 65494 172454 100938
rect 181794 111454 182414 146898
rect 189234 154894 189854 190338
rect 192954 194614 193574 230058
rect 196674 234334 197294 269778
rect 204114 277774 204734 313218
rect 207834 317494 208454 352938
rect 217794 363454 218414 398898
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221008 378334 221328 378366
rect 221008 378098 221050 378334
rect 221286 378098 221328 378334
rect 221008 378014 221328 378098
rect 221008 377778 221050 378014
rect 221286 377778 221328 378014
rect 221008 377746 221328 377778
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 215888 338614 216208 338646
rect 215888 338378 215930 338614
rect 216166 338378 216208 338614
rect 215888 338294 216208 338378
rect 215888 338058 215930 338294
rect 216166 338058 216208 338294
rect 215888 338026 216208 338058
rect 210768 334894 211088 334926
rect 210768 334658 210810 334894
rect 211046 334658 211088 334894
rect 210768 334574 211088 334658
rect 210768 334338 210810 334574
rect 211046 334338 211088 334574
rect 210768 334306 211088 334338
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 205648 295174 205968 295206
rect 205648 294938 205690 295174
rect 205926 294938 205968 295174
rect 205648 294854 205968 294938
rect 205648 294618 205690 294854
rect 205926 294618 205968 294854
rect 205648 294586 205968 294618
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 200528 255454 200848 255486
rect 200528 255218 200570 255454
rect 200806 255218 200848 255454
rect 200528 255134 200848 255218
rect 200528 254898 200570 255134
rect 200806 254898 200848 255134
rect 200528 254866 200848 254898
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 195408 202054 195728 202086
rect 195408 201818 195450 202054
rect 195686 201818 195728 202054
rect 195408 201734 195728 201818
rect 195408 201498 195450 201734
rect 195686 201498 195728 201734
rect 195408 201466 195728 201498
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 190288 162334 190608 162366
rect 190288 162098 190330 162334
rect 190566 162098 190608 162334
rect 190288 162014 190608 162098
rect 190288 161778 190330 162014
rect 190566 161778 190608 162014
rect 190288 161746 190608 161778
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 185168 122614 185488 122646
rect 185168 122378 185210 122614
rect 185446 122378 185488 122614
rect 185168 122294 185488 122378
rect 185168 122058 185210 122294
rect 185446 122058 185488 122294
rect 185168 122026 185488 122058
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 180048 82894 180368 82926
rect 180048 82658 180090 82894
rect 180326 82658 180368 82894
rect 180048 82574 180368 82658
rect 180048 82338 180090 82574
rect 180326 82338 180368 82574
rect 180048 82306 180368 82338
rect 174928 79174 175248 79206
rect 174928 78938 174970 79174
rect 175206 78938 175248 79174
rect 174928 78854 175248 78938
rect 174928 78618 174970 78854
rect 175206 78618 175248 78854
rect 174928 78586 175248 78618
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 169808 39454 170128 39486
rect 169808 39218 169850 39454
rect 170086 39218 170128 39454
rect 169808 39134 170128 39218
rect 169808 38898 169850 39134
rect 170086 38898 170128 39134
rect 169808 38866 170128 38898
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 164688 22054 165008 22086
rect 164688 21818 164730 22054
rect 164966 21818 165008 22054
rect 164688 21734 165008 21818
rect 164688 21498 164730 21734
rect 164966 21498 165008 21734
rect 164688 21466 165008 21498
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 -1306 150134 2988
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 -5146 165014 2988
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 64938
rect 181794 75454 182414 110898
rect 189234 118894 189854 154338
rect 192954 158614 193574 194058
rect 196674 198334 197294 233778
rect 204114 241774 204734 277218
rect 207834 281494 208454 316938
rect 217794 327454 218414 362898
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221008 342334 221328 342366
rect 221008 342098 221050 342334
rect 221286 342098 221328 342334
rect 221008 342014 221328 342098
rect 221008 341778 221050 342014
rect 221286 341778 221328 342014
rect 221008 341746 221328 341778
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 215888 302614 216208 302646
rect 215888 302378 215930 302614
rect 216166 302378 216208 302614
rect 215888 302294 216208 302378
rect 215888 302058 215930 302294
rect 216166 302058 216208 302294
rect 215888 302026 216208 302058
rect 210768 298894 211088 298926
rect 210768 298658 210810 298894
rect 211046 298658 211088 298894
rect 210768 298574 211088 298658
rect 210768 298338 210810 298574
rect 211046 298338 211088 298574
rect 210768 298306 211088 298338
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 205648 259174 205968 259206
rect 205648 258938 205690 259174
rect 205926 258938 205968 259174
rect 205648 258854 205968 258938
rect 205648 258618 205690 258854
rect 205926 258618 205968 258854
rect 205648 258586 205968 258618
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 200528 219454 200848 219486
rect 200528 219218 200570 219454
rect 200806 219218 200848 219454
rect 200528 219134 200848 219218
rect 200528 218898 200570 219134
rect 200806 218898 200848 219134
rect 200528 218866 200848 218898
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 195408 166054 195728 166086
rect 195408 165818 195450 166054
rect 195686 165818 195728 166054
rect 195408 165734 195728 165818
rect 195408 165498 195450 165734
rect 195686 165498 195728 165734
rect 195408 165466 195728 165498
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 190288 126334 190608 126366
rect 190288 126098 190330 126334
rect 190566 126098 190608 126334
rect 190288 126014 190608 126098
rect 190288 125778 190330 126014
rect 190566 125778 190608 126014
rect 190288 125746 190608 125778
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 185168 86614 185488 86646
rect 185168 86378 185210 86614
rect 185446 86378 185488 86614
rect 185168 86294 185488 86378
rect 185168 86058 185210 86294
rect 185446 86058 185488 86294
rect 185168 86026 185488 86058
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 180048 46894 180368 46926
rect 180048 46658 180090 46894
rect 180326 46658 180368 46894
rect 180048 46574 180368 46658
rect 180048 46338 180090 46574
rect 180326 46338 180368 46574
rect 180048 46306 180368 46338
rect 174928 43174 175248 43206
rect 174928 42938 174970 43174
rect 175206 42938 175248 43174
rect 174928 42854 175248 42938
rect 174928 42618 174970 42854
rect 175206 42618 175248 42854
rect 174928 42586 175248 42618
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 181794 39454 182414 74898
rect 189234 82894 189854 118338
rect 192954 122614 193574 158058
rect 196674 162334 197294 197778
rect 204114 205774 204734 241218
rect 207834 245494 208454 280938
rect 217794 291454 218414 326898
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221008 306334 221328 306366
rect 221008 306098 221050 306334
rect 221286 306098 221328 306334
rect 221008 306014 221328 306098
rect 221008 305778 221050 306014
rect 221286 305778 221328 306014
rect 221008 305746 221328 305778
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 215888 266614 216208 266646
rect 215888 266378 215930 266614
rect 216166 266378 216208 266614
rect 215888 266294 216208 266378
rect 215888 266058 215930 266294
rect 216166 266058 216208 266294
rect 215888 266026 216208 266058
rect 210768 262894 211088 262926
rect 210768 262658 210810 262894
rect 211046 262658 211088 262894
rect 210768 262574 211088 262658
rect 210768 262338 210810 262574
rect 211046 262338 211088 262574
rect 210768 262306 211088 262338
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 205648 223174 205968 223206
rect 205648 222938 205690 223174
rect 205926 222938 205968 223174
rect 205648 222854 205968 222938
rect 205648 222618 205690 222854
rect 205926 222618 205968 222854
rect 205648 222586 205968 222618
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 200528 183454 200848 183486
rect 200528 183218 200570 183454
rect 200806 183218 200848 183454
rect 200528 183134 200848 183218
rect 200528 182898 200570 183134
rect 200806 182898 200848 183134
rect 200528 182866 200848 182898
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 195408 130054 195728 130086
rect 195408 129818 195450 130054
rect 195686 129818 195728 130054
rect 195408 129734 195728 129818
rect 195408 129498 195450 129734
rect 195686 129498 195728 129734
rect 195408 129466 195728 129498
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 190288 90334 190608 90366
rect 190288 90098 190330 90334
rect 190566 90098 190608 90334
rect 190288 90014 190608 90098
rect 190288 89778 190330 90014
rect 190566 89778 190608 90014
rect 190288 89746 190608 89778
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 185168 50614 185488 50646
rect 185168 50378 185210 50614
rect 185446 50378 185488 50614
rect 185168 50294 185488 50378
rect 185168 50058 185210 50294
rect 185446 50058 185488 50294
rect 185168 50026 185488 50058
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 180048 10894 180368 10926
rect 180048 10658 180090 10894
rect 180326 10658 180368 10894
rect 180048 10574 180368 10658
rect 180048 10338 180090 10574
rect 180326 10338 180368 10574
rect 180048 10306 180368 10338
rect 174928 7174 175248 7206
rect 174928 6938 174970 7174
rect 175206 6938 175248 7174
rect 174928 6854 175248 6938
rect 174928 6618 174970 6854
rect 175206 6618 175248 6854
rect 174928 6586 175248 6618
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 3454 182414 38898
rect 189234 46894 189854 82338
rect 192954 86614 193574 122058
rect 196674 126334 197294 161778
rect 204114 169774 204734 205218
rect 207834 209494 208454 244938
rect 217794 255454 218414 290898
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221008 270334 221328 270366
rect 221008 270098 221050 270334
rect 221286 270098 221328 270334
rect 221008 270014 221328 270098
rect 221008 269778 221050 270014
rect 221286 269778 221328 270014
rect 221008 269746 221328 269778
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 215888 230614 216208 230646
rect 215888 230378 215930 230614
rect 216166 230378 216208 230614
rect 215888 230294 216208 230378
rect 215888 230058 215930 230294
rect 216166 230058 216208 230294
rect 215888 230026 216208 230058
rect 210768 226894 211088 226926
rect 210768 226658 210810 226894
rect 211046 226658 211088 226894
rect 210768 226574 211088 226658
rect 210768 226338 210810 226574
rect 211046 226338 211088 226574
rect 210768 226306 211088 226338
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 205648 187174 205968 187206
rect 205648 186938 205690 187174
rect 205926 186938 205968 187174
rect 205648 186854 205968 186938
rect 205648 186618 205690 186854
rect 205926 186618 205968 186854
rect 205648 186586 205968 186618
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 200528 147454 200848 147486
rect 200528 147218 200570 147454
rect 200806 147218 200848 147454
rect 200528 147134 200848 147218
rect 200528 146898 200570 147134
rect 200806 146898 200848 147134
rect 200528 146866 200848 146898
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 195408 94054 195728 94086
rect 195408 93818 195450 94054
rect 195686 93818 195728 94054
rect 195408 93734 195728 93818
rect 195408 93498 195450 93734
rect 195686 93498 195728 93734
rect 195408 93466 195728 93498
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 190288 54334 190608 54366
rect 190288 54098 190330 54334
rect 190566 54098 190608 54334
rect 190288 54014 190608 54098
rect 190288 53778 190330 54014
rect 190566 53778 190608 54014
rect 190288 53746 190608 53778
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 185168 14614 185488 14646
rect 185168 14378 185210 14614
rect 185446 14378 185488 14614
rect 185168 14294 185488 14378
rect 185168 14058 185210 14294
rect 185446 14058 185488 14294
rect 185168 14026 185488 14058
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 189234 10894 189854 46338
rect 192954 50614 193574 86058
rect 196674 90334 197294 125778
rect 204114 133774 204734 169218
rect 207834 173494 208454 208938
rect 217794 219454 218414 254898
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221008 234334 221328 234366
rect 221008 234098 221050 234334
rect 221286 234098 221328 234334
rect 221008 234014 221328 234098
rect 221008 233778 221050 234014
rect 221286 233778 221328 234014
rect 221008 233746 221328 233778
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 215888 194614 216208 194646
rect 215888 194378 215930 194614
rect 216166 194378 216208 194614
rect 215888 194294 216208 194378
rect 215888 194058 215930 194294
rect 216166 194058 216208 194294
rect 215888 194026 216208 194058
rect 210768 190894 211088 190926
rect 210768 190658 210810 190894
rect 211046 190658 211088 190894
rect 210768 190574 211088 190658
rect 210768 190338 210810 190574
rect 211046 190338 211088 190574
rect 210768 190306 211088 190338
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 205648 151174 205968 151206
rect 205648 150938 205690 151174
rect 205926 150938 205968 151174
rect 205648 150854 205968 150938
rect 205648 150618 205690 150854
rect 205926 150618 205968 150854
rect 205648 150586 205968 150618
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 200528 111454 200848 111486
rect 200528 111218 200570 111454
rect 200806 111218 200848 111454
rect 200528 111134 200848 111218
rect 200528 110898 200570 111134
rect 200806 110898 200848 111134
rect 200528 110866 200848 110898
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 195408 58054 195728 58086
rect 195408 57818 195450 58054
rect 195686 57818 195728 58054
rect 195408 57734 195728 57818
rect 195408 57498 195450 57734
rect 195686 57498 195728 57734
rect 195408 57466 195728 57498
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 190288 18334 190608 18366
rect 190288 18098 190330 18334
rect 190566 18098 190608 18334
rect 190288 18014 190608 18098
rect 190288 17778 190330 18014
rect 190566 17778 190608 18014
rect 190288 17746 190608 17778
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 -1306 186134 2988
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 50058
rect 196674 54334 197294 89778
rect 204114 97774 204734 133218
rect 207834 137494 208454 172938
rect 217794 183454 218414 218898
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221008 198334 221328 198366
rect 221008 198098 221050 198334
rect 221286 198098 221328 198334
rect 221008 198014 221328 198098
rect 221008 197778 221050 198014
rect 221286 197778 221328 198014
rect 221008 197746 221328 197778
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 215888 158614 216208 158646
rect 215888 158378 215930 158614
rect 216166 158378 216208 158614
rect 215888 158294 216208 158378
rect 215888 158058 215930 158294
rect 216166 158058 216208 158294
rect 215888 158026 216208 158058
rect 210768 154894 211088 154926
rect 210768 154658 210810 154894
rect 211046 154658 211088 154894
rect 210768 154574 211088 154658
rect 210768 154338 210810 154574
rect 211046 154338 211088 154574
rect 210768 154306 211088 154338
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 205648 115174 205968 115206
rect 205648 114938 205690 115174
rect 205926 114938 205968 115174
rect 205648 114854 205968 114938
rect 205648 114618 205690 114854
rect 205926 114618 205968 114854
rect 205648 114586 205968 114618
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 200528 75454 200848 75486
rect 200528 75218 200570 75454
rect 200806 75218 200848 75454
rect 200528 75134 200848 75218
rect 200528 74898 200570 75134
rect 200806 74898 200848 75134
rect 200528 74866 200848 74898
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 195408 22054 195728 22086
rect 195408 21818 195450 22054
rect 195686 21818 195728 22054
rect 195408 21734 195728 21818
rect 195408 21498 195450 21734
rect 195686 21498 195728 21734
rect 195408 21466 195728 21498
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 53778
rect 204114 61774 204734 97218
rect 207834 101494 208454 136938
rect 217794 147454 218414 182898
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221008 162334 221328 162366
rect 221008 162098 221050 162334
rect 221286 162098 221328 162334
rect 221008 162014 221328 162098
rect 221008 161778 221050 162014
rect 221286 161778 221328 162014
rect 221008 161746 221328 161778
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 215888 122614 216208 122646
rect 215888 122378 215930 122614
rect 216166 122378 216208 122614
rect 215888 122294 216208 122378
rect 215888 122058 215930 122294
rect 216166 122058 216208 122294
rect 215888 122026 216208 122058
rect 210768 118894 211088 118926
rect 210768 118658 210810 118894
rect 211046 118658 211088 118894
rect 210768 118574 211088 118658
rect 210768 118338 210810 118574
rect 211046 118338 211088 118574
rect 210768 118306 211088 118338
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 205648 79174 205968 79206
rect 205648 78938 205690 79174
rect 205926 78938 205968 79174
rect 205648 78854 205968 78938
rect 205648 78618 205690 78854
rect 205926 78618 205968 78854
rect 205648 78586 205968 78618
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 200528 39454 200848 39486
rect 200528 39218 200570 39454
rect 200806 39218 200848 39454
rect 200528 39134 200848 39218
rect 200528 38898 200570 39134
rect 200806 38898 200848 39134
rect 200528 38866 200848 38898
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 204114 25774 204734 61218
rect 207834 65494 208454 100938
rect 217794 111454 218414 146898
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221008 126334 221328 126366
rect 221008 126098 221050 126334
rect 221286 126098 221328 126334
rect 221008 126014 221328 126098
rect 221008 125778 221050 126014
rect 221286 125778 221328 126014
rect 221008 125746 221328 125778
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 215888 86614 216208 86646
rect 215888 86378 215930 86614
rect 216166 86378 216208 86614
rect 215888 86294 216208 86378
rect 215888 86058 215930 86294
rect 216166 86058 216208 86294
rect 215888 86026 216208 86058
rect 210768 82894 211088 82926
rect 210768 82658 210810 82894
rect 211046 82658 211088 82894
rect 210768 82574 211088 82658
rect 210768 82338 210810 82574
rect 211046 82338 211088 82574
rect 210768 82306 211088 82338
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 205648 43174 205968 43206
rect 205648 42938 205690 43174
rect 205926 42938 205968 43174
rect 205648 42854 205968 42938
rect 205648 42618 205690 42854
rect 205926 42618 205968 42854
rect 205648 42586 205968 42618
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 -5146 201014 2988
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 -6106 204734 25218
rect 207834 29494 208454 64938
rect 217794 75454 218414 110898
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221008 90334 221328 90366
rect 221008 90098 221050 90334
rect 221286 90098 221328 90334
rect 221008 90014 221328 90098
rect 221008 89778 221050 90014
rect 221286 89778 221328 90014
rect 221008 89746 221328 89778
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 215888 50614 216208 50646
rect 215888 50378 215930 50614
rect 216166 50378 216208 50614
rect 215888 50294 216208 50378
rect 215888 50058 215930 50294
rect 216166 50058 216208 50294
rect 215888 50026 216208 50058
rect 210768 46894 211088 46926
rect 210768 46658 210810 46894
rect 211046 46658 211088 46894
rect 210768 46574 211088 46658
rect 210768 46338 210810 46574
rect 211046 46338 211088 46574
rect 210768 46306 211088 46338
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 205648 7174 205968 7206
rect 205648 6938 205690 7174
rect 205926 6938 205968 7174
rect 205648 6854 205968 6938
rect 205648 6618 205690 6854
rect 205926 6618 205968 6854
rect 205648 6586 205968 6618
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 -7066 208454 28938
rect 217794 39454 218414 74898
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221008 54334 221328 54366
rect 221008 54098 221050 54334
rect 221286 54098 221328 54334
rect 221008 54014 221328 54098
rect 221008 53778 221050 54014
rect 221286 53778 221328 54014
rect 221008 53746 221328 53778
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 215888 14614 216208 14646
rect 215888 14378 215930 14614
rect 216166 14378 216208 14614
rect 215888 14294 216208 14378
rect 215888 14058 215930 14294
rect 216166 14058 216208 14294
rect 215888 14026 216208 14058
rect 210768 10894 211088 10926
rect 210768 10658 210810 10894
rect 211046 10658 211088 10894
rect 210768 10574 211088 10658
rect 210768 10338 210810 10574
rect 211046 10338 211088 10574
rect 210768 10306 211088 10338
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 3454 218414 38898
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221008 18334 221328 18366
rect 221008 18098 221050 18334
rect 221286 18098 221328 18334
rect 221008 18014 221328 18098
rect 221008 17778 221050 18014
rect 221286 17778 221328 18014
rect 221008 17746 221328 17778
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 226128 598054 226448 598086
rect 226128 597818 226170 598054
rect 226406 597818 226448 598054
rect 226128 597734 226448 597818
rect 226128 597498 226170 597734
rect 226406 597498 226448 597734
rect 226128 597466 226448 597498
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 226128 562054 226448 562086
rect 226128 561818 226170 562054
rect 226406 561818 226448 562054
rect 226128 561734 226448 561818
rect 226128 561498 226170 561734
rect 226406 561498 226448 561734
rect 226128 561466 226448 561498
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 228954 554614 229574 590058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 594334 233294 629778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 602500 237014 633498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 232674 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 233294 594334
rect 232674 594014 233294 594098
rect 232674 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 233294 594014
rect 231248 579454 231568 579486
rect 231248 579218 231290 579454
rect 231526 579218 231568 579454
rect 231248 579134 231568 579218
rect 231248 578898 231290 579134
rect 231526 578898 231568 579134
rect 231248 578866 231568 578898
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 226128 526054 226448 526086
rect 226128 525818 226170 526054
rect 226406 525818 226448 526054
rect 226128 525734 226448 525818
rect 226128 525498 226170 525734
rect 226406 525498 226448 525734
rect 226128 525466 226448 525498
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 228954 518614 229574 554058
rect 232674 558334 233294 593778
rect 240114 601774 240734 637218
rect 240114 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 240734 601774
rect 240114 601454 240734 601538
rect 240114 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 240734 601454
rect 236368 583174 236688 583206
rect 236368 582938 236410 583174
rect 236646 582938 236688 583174
rect 236368 582854 236688 582938
rect 236368 582618 236410 582854
rect 236646 582618 236688 582854
rect 236368 582586 236688 582618
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 231248 543454 231568 543486
rect 231248 543218 231290 543454
rect 231526 543218 231568 543454
rect 231248 543134 231568 543218
rect 231248 542898 231290 543134
rect 231526 542898 231568 543134
rect 231248 542866 231568 542898
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 226128 490054 226448 490086
rect 226128 489818 226170 490054
rect 226406 489818 226448 490054
rect 226128 489734 226448 489818
rect 226128 489498 226170 489734
rect 226406 489498 226448 489734
rect 226128 489466 226448 489498
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 228954 482614 229574 518058
rect 232674 522334 233294 557778
rect 240114 565774 240734 601218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 605494 244454 640938
rect 243834 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 244454 605494
rect 243834 605174 244454 605258
rect 243834 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 244454 605174
rect 241488 586894 241808 586926
rect 241488 586658 241530 586894
rect 241766 586658 241808 586894
rect 241488 586574 241808 586658
rect 241488 586338 241530 586574
rect 241766 586338 241808 586574
rect 241488 586306 241808 586338
rect 240114 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 240734 565774
rect 240114 565454 240734 565538
rect 240114 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 240734 565454
rect 236368 547174 236688 547206
rect 236368 546938 236410 547174
rect 236646 546938 236688 547174
rect 236368 546854 236688 546938
rect 236368 546618 236410 546854
rect 236646 546618 236688 546854
rect 236368 546586 236688 546618
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 231248 507454 231568 507486
rect 231248 507218 231290 507454
rect 231526 507218 231568 507454
rect 231248 507134 231568 507218
rect 231248 506898 231290 507134
rect 231526 506898 231568 507134
rect 231248 506866 231568 506898
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 226128 454054 226448 454086
rect 226128 453818 226170 454054
rect 226406 453818 226448 454054
rect 226128 453734 226448 453818
rect 226128 453498 226170 453734
rect 226406 453498 226448 453734
rect 226128 453466 226448 453498
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 228954 446614 229574 482058
rect 232674 486334 233294 521778
rect 240114 529774 240734 565218
rect 243834 569494 244454 604938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 251728 594334 252048 594366
rect 251728 594098 251770 594334
rect 252006 594098 252048 594334
rect 251728 594014 252048 594098
rect 251728 593778 251770 594014
rect 252006 593778 252048 594014
rect 251728 593746 252048 593778
rect 246608 590614 246928 590646
rect 246608 590378 246650 590614
rect 246886 590378 246928 590614
rect 246608 590294 246928 590378
rect 246608 590058 246650 590294
rect 246886 590058 246928 590294
rect 246608 590026 246928 590058
rect 243834 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 244454 569494
rect 243834 569174 244454 569258
rect 243834 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 244454 569174
rect 241488 550894 241808 550926
rect 241488 550658 241530 550894
rect 241766 550658 241808 550894
rect 241488 550574 241808 550658
rect 241488 550338 241530 550574
rect 241766 550338 241808 550574
rect 241488 550306 241808 550338
rect 240114 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 240734 529774
rect 240114 529454 240734 529538
rect 240114 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 240734 529454
rect 236368 511174 236688 511206
rect 236368 510938 236410 511174
rect 236646 510938 236688 511174
rect 236368 510854 236688 510938
rect 236368 510618 236410 510854
rect 236646 510618 236688 510854
rect 236368 510586 236688 510618
rect 232674 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 233294 486334
rect 232674 486014 233294 486098
rect 232674 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 233294 486014
rect 231248 471454 231568 471486
rect 231248 471218 231290 471454
rect 231526 471218 231568 471454
rect 231248 471134 231568 471218
rect 231248 470898 231290 471134
rect 231526 470898 231568 471134
rect 231248 470866 231568 470898
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 226128 418054 226448 418086
rect 226128 417818 226170 418054
rect 226406 417818 226448 418054
rect 226128 417734 226448 417818
rect 226128 417498 226170 417734
rect 226406 417498 226448 417734
rect 226128 417466 226448 417498
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 228954 410614 229574 446058
rect 232674 450334 233294 485778
rect 240114 493774 240734 529218
rect 243834 533494 244454 568938
rect 253794 579454 254414 614898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 256848 598054 257168 598086
rect 256848 597818 256890 598054
rect 257126 597818 257168 598054
rect 256848 597734 257168 597818
rect 256848 597498 256890 597734
rect 257126 597498 257168 597734
rect 256848 597466 257168 597498
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 251728 558334 252048 558366
rect 251728 558098 251770 558334
rect 252006 558098 252048 558334
rect 251728 558014 252048 558098
rect 251728 557778 251770 558014
rect 252006 557778 252048 558014
rect 251728 557746 252048 557778
rect 246608 554614 246928 554646
rect 246608 554378 246650 554614
rect 246886 554378 246928 554614
rect 246608 554294 246928 554378
rect 246608 554058 246650 554294
rect 246886 554058 246928 554294
rect 246608 554026 246928 554058
rect 243834 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 244454 533494
rect 243834 533174 244454 533258
rect 243834 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 244454 533174
rect 241488 514894 241808 514926
rect 241488 514658 241530 514894
rect 241766 514658 241808 514894
rect 241488 514574 241808 514658
rect 241488 514338 241530 514574
rect 241766 514338 241808 514574
rect 241488 514306 241808 514338
rect 240114 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 240734 493774
rect 240114 493454 240734 493538
rect 240114 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 240734 493454
rect 236368 475174 236688 475206
rect 236368 474938 236410 475174
rect 236646 474938 236688 475174
rect 236368 474854 236688 474938
rect 236368 474618 236410 474854
rect 236646 474618 236688 474854
rect 236368 474586 236688 474618
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 231248 435454 231568 435486
rect 231248 435218 231290 435454
rect 231526 435218 231568 435454
rect 231248 435134 231568 435218
rect 231248 434898 231290 435134
rect 231526 434898 231568 435134
rect 231248 434866 231568 434898
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 226128 382054 226448 382086
rect 226128 381818 226170 382054
rect 226406 381818 226448 382054
rect 226128 381734 226448 381818
rect 226128 381498 226170 381734
rect 226406 381498 226448 381734
rect 226128 381466 226448 381498
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 228954 374614 229574 410058
rect 232674 414334 233294 449778
rect 240114 457774 240734 493218
rect 243834 497494 244454 532938
rect 253794 543454 254414 578898
rect 257514 583174 258134 618618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 602500 261854 622338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 256848 562054 257168 562086
rect 256848 561818 256890 562054
rect 257126 561818 257168 562054
rect 256848 561734 257168 561818
rect 256848 561498 256890 561734
rect 257126 561498 257168 561734
rect 256848 561466 257168 561498
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 251728 522334 252048 522366
rect 251728 522098 251770 522334
rect 252006 522098 252048 522334
rect 251728 522014 252048 522098
rect 251728 521778 251770 522014
rect 252006 521778 252048 522014
rect 251728 521746 252048 521778
rect 246608 518614 246928 518646
rect 246608 518378 246650 518614
rect 246886 518378 246928 518614
rect 246608 518294 246928 518378
rect 246608 518058 246650 518294
rect 246886 518058 246928 518294
rect 246608 518026 246928 518058
rect 243834 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 244454 497494
rect 243834 497174 244454 497258
rect 243834 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 244454 497174
rect 241488 478894 241808 478926
rect 241488 478658 241530 478894
rect 241766 478658 241808 478894
rect 241488 478574 241808 478658
rect 241488 478338 241530 478574
rect 241766 478338 241808 478574
rect 241488 478306 241808 478338
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 236368 439174 236688 439206
rect 236368 438938 236410 439174
rect 236646 438938 236688 439174
rect 236368 438854 236688 438938
rect 236368 438618 236410 438854
rect 236646 438618 236688 438854
rect 236368 438586 236688 438618
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 231248 399454 231568 399486
rect 231248 399218 231290 399454
rect 231526 399218 231568 399454
rect 231248 399134 231568 399218
rect 231248 398898 231290 399134
rect 231526 398898 231568 399134
rect 231248 398866 231568 398898
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 226128 346054 226448 346086
rect 226128 345818 226170 346054
rect 226406 345818 226448 346054
rect 226128 345734 226448 345818
rect 226128 345498 226170 345734
rect 226406 345498 226448 345734
rect 226128 345466 226448 345498
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 228954 338614 229574 374058
rect 232674 378334 233294 413778
rect 240114 421774 240734 457218
rect 243834 461494 244454 496938
rect 253794 507454 254414 542898
rect 257514 547174 258134 582618
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 261968 579454 262288 579486
rect 261968 579218 262010 579454
rect 262246 579218 262288 579454
rect 261968 579134 262288 579218
rect 261968 578898 262010 579134
rect 262246 578898 262288 579134
rect 261968 578866 262288 578898
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 256848 526054 257168 526086
rect 256848 525818 256890 526054
rect 257126 525818 257168 526054
rect 256848 525734 257168 525818
rect 256848 525498 256890 525734
rect 257126 525498 257168 525734
rect 256848 525466 257168 525498
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 251728 486334 252048 486366
rect 251728 486098 251770 486334
rect 252006 486098 252048 486334
rect 251728 486014 252048 486098
rect 251728 485778 251770 486014
rect 252006 485778 252048 486014
rect 251728 485746 252048 485778
rect 246608 482614 246928 482646
rect 246608 482378 246650 482614
rect 246886 482378 246928 482614
rect 246608 482294 246928 482378
rect 246608 482058 246650 482294
rect 246886 482058 246928 482294
rect 246608 482026 246928 482058
rect 243834 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 244454 461494
rect 243834 461174 244454 461258
rect 243834 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 244454 461174
rect 241488 442894 241808 442926
rect 241488 442658 241530 442894
rect 241766 442658 241808 442894
rect 241488 442574 241808 442658
rect 241488 442338 241530 442574
rect 241766 442338 241808 442574
rect 241488 442306 241808 442338
rect 240114 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 240734 421774
rect 240114 421454 240734 421538
rect 240114 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 240734 421454
rect 236368 403174 236688 403206
rect 236368 402938 236410 403174
rect 236646 402938 236688 403174
rect 236368 402854 236688 402938
rect 236368 402618 236410 402854
rect 236646 402618 236688 402854
rect 236368 402586 236688 402618
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 231248 363454 231568 363486
rect 231248 363218 231290 363454
rect 231526 363218 231568 363454
rect 231248 363134 231568 363218
rect 231248 362898 231290 363134
rect 231526 362898 231568 363134
rect 231248 362866 231568 362898
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 226128 310054 226448 310086
rect 226128 309818 226170 310054
rect 226406 309818 226448 310054
rect 226128 309734 226448 309818
rect 226128 309498 226170 309734
rect 226406 309498 226448 309734
rect 226128 309466 226448 309498
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 228954 302614 229574 338058
rect 232674 342334 233294 377778
rect 240114 385774 240734 421218
rect 243834 425494 244454 460938
rect 253794 471454 254414 506898
rect 257514 511174 258134 546618
rect 264954 554614 265574 590058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 268674 594334 269294 629778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 272394 602500 273014 633498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 268674 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 269294 594334
rect 268674 594014 269294 594098
rect 268674 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 269294 594014
rect 267088 583174 267408 583206
rect 267088 582938 267130 583174
rect 267366 582938 267408 583174
rect 267088 582854 267408 582938
rect 267088 582618 267130 582854
rect 267366 582618 267408 582854
rect 267088 582586 267408 582618
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 261968 543454 262288 543486
rect 261968 543218 262010 543454
rect 262246 543218 262288 543454
rect 261968 543134 262288 543218
rect 261968 542898 262010 543134
rect 262246 542898 262288 543134
rect 261968 542866 262288 542898
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 256848 490054 257168 490086
rect 256848 489818 256890 490054
rect 257126 489818 257168 490054
rect 256848 489734 257168 489818
rect 256848 489498 256890 489734
rect 257126 489498 257168 489734
rect 256848 489466 257168 489498
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 251728 450334 252048 450366
rect 251728 450098 251770 450334
rect 252006 450098 252048 450334
rect 251728 450014 252048 450098
rect 251728 449778 251770 450014
rect 252006 449778 252048 450014
rect 251728 449746 252048 449778
rect 246608 446614 246928 446646
rect 246608 446378 246650 446614
rect 246886 446378 246928 446614
rect 246608 446294 246928 446378
rect 246608 446058 246650 446294
rect 246886 446058 246928 446294
rect 246608 446026 246928 446058
rect 243834 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 244454 425494
rect 243834 425174 244454 425258
rect 243834 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 244454 425174
rect 241488 406894 241808 406926
rect 241488 406658 241530 406894
rect 241766 406658 241808 406894
rect 241488 406574 241808 406658
rect 241488 406338 241530 406574
rect 241766 406338 241808 406574
rect 241488 406306 241808 406338
rect 240114 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 240734 385774
rect 240114 385454 240734 385538
rect 240114 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 240734 385454
rect 236368 367174 236688 367206
rect 236368 366938 236410 367174
rect 236646 366938 236688 367174
rect 236368 366854 236688 366938
rect 236368 366618 236410 366854
rect 236646 366618 236688 366854
rect 236368 366586 236688 366618
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 231248 327454 231568 327486
rect 231248 327218 231290 327454
rect 231526 327218 231568 327454
rect 231248 327134 231568 327218
rect 231248 326898 231290 327134
rect 231526 326898 231568 327134
rect 231248 326866 231568 326898
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 226128 274054 226448 274086
rect 226128 273818 226170 274054
rect 226406 273818 226448 274054
rect 226128 273734 226448 273818
rect 226128 273498 226170 273734
rect 226406 273498 226448 273734
rect 226128 273466 226448 273498
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 228954 266614 229574 302058
rect 232674 306334 233294 341778
rect 240114 349774 240734 385218
rect 243834 389494 244454 424938
rect 253794 435454 254414 470898
rect 257514 475174 258134 510618
rect 264954 518614 265574 554058
rect 268674 558334 269294 593778
rect 276114 601774 276734 637218
rect 276114 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 276734 601774
rect 276114 601454 276734 601538
rect 276114 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 276734 601454
rect 272208 586894 272528 586926
rect 272208 586658 272250 586894
rect 272486 586658 272528 586894
rect 272208 586574 272528 586658
rect 272208 586338 272250 586574
rect 272486 586338 272528 586574
rect 272208 586306 272528 586338
rect 268674 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 269294 558334
rect 268674 558014 269294 558098
rect 268674 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 269294 558014
rect 267088 547174 267408 547206
rect 267088 546938 267130 547174
rect 267366 546938 267408 547174
rect 267088 546854 267408 546938
rect 267088 546618 267130 546854
rect 267366 546618 267408 546854
rect 267088 546586 267408 546618
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 261968 507454 262288 507486
rect 261968 507218 262010 507454
rect 262246 507218 262288 507454
rect 261968 507134 262288 507218
rect 261968 506898 262010 507134
rect 262246 506898 262288 507134
rect 261968 506866 262288 506898
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 256848 454054 257168 454086
rect 256848 453818 256890 454054
rect 257126 453818 257168 454054
rect 256848 453734 257168 453818
rect 256848 453498 256890 453734
rect 257126 453498 257168 453734
rect 256848 453466 257168 453498
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 251728 414334 252048 414366
rect 251728 414098 251770 414334
rect 252006 414098 252048 414334
rect 251728 414014 252048 414098
rect 251728 413778 251770 414014
rect 252006 413778 252048 414014
rect 251728 413746 252048 413778
rect 246608 410614 246928 410646
rect 246608 410378 246650 410614
rect 246886 410378 246928 410614
rect 246608 410294 246928 410378
rect 246608 410058 246650 410294
rect 246886 410058 246928 410294
rect 246608 410026 246928 410058
rect 243834 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 244454 389494
rect 243834 389174 244454 389258
rect 243834 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 244454 389174
rect 241488 370894 241808 370926
rect 241488 370658 241530 370894
rect 241766 370658 241808 370894
rect 241488 370574 241808 370658
rect 241488 370338 241530 370574
rect 241766 370338 241808 370574
rect 241488 370306 241808 370338
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 236368 331174 236688 331206
rect 236368 330938 236410 331174
rect 236646 330938 236688 331174
rect 236368 330854 236688 330938
rect 236368 330618 236410 330854
rect 236646 330618 236688 330854
rect 236368 330586 236688 330618
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 231248 291454 231568 291486
rect 231248 291218 231290 291454
rect 231526 291218 231568 291454
rect 231248 291134 231568 291218
rect 231248 290898 231290 291134
rect 231526 290898 231568 291134
rect 231248 290866 231568 290898
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 226128 238054 226448 238086
rect 226128 237818 226170 238054
rect 226406 237818 226448 238054
rect 226128 237734 226448 237818
rect 226128 237498 226170 237734
rect 226406 237498 226448 237734
rect 226128 237466 226448 237498
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 228954 230614 229574 266058
rect 232674 270334 233294 305778
rect 240114 313774 240734 349218
rect 243834 353494 244454 388938
rect 253794 399454 254414 434898
rect 257514 439174 258134 474618
rect 264954 482614 265574 518058
rect 268674 522334 269294 557778
rect 276114 565774 276734 601218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 605494 280454 640938
rect 279834 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 280454 605494
rect 279834 605174 280454 605258
rect 279834 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 280454 605174
rect 277328 590614 277648 590646
rect 277328 590378 277370 590614
rect 277606 590378 277648 590614
rect 277328 590294 277648 590378
rect 277328 590058 277370 590294
rect 277606 590058 277648 590294
rect 277328 590026 277648 590058
rect 276114 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 276734 565774
rect 276114 565454 276734 565538
rect 276114 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 276734 565454
rect 272208 550894 272528 550926
rect 272208 550658 272250 550894
rect 272486 550658 272528 550894
rect 272208 550574 272528 550658
rect 272208 550338 272250 550574
rect 272486 550338 272528 550574
rect 272208 550306 272528 550338
rect 268674 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 269294 522334
rect 268674 522014 269294 522098
rect 268674 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 269294 522014
rect 267088 511174 267408 511206
rect 267088 510938 267130 511174
rect 267366 510938 267408 511174
rect 267088 510854 267408 510938
rect 267088 510618 267130 510854
rect 267366 510618 267408 510854
rect 267088 510586 267408 510618
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 261968 471454 262288 471486
rect 261968 471218 262010 471454
rect 262246 471218 262288 471454
rect 261968 471134 262288 471218
rect 261968 470898 262010 471134
rect 262246 470898 262288 471134
rect 261968 470866 262288 470898
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 256848 418054 257168 418086
rect 256848 417818 256890 418054
rect 257126 417818 257168 418054
rect 256848 417734 257168 417818
rect 256848 417498 256890 417734
rect 257126 417498 257168 417734
rect 256848 417466 257168 417498
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 251728 378334 252048 378366
rect 251728 378098 251770 378334
rect 252006 378098 252048 378334
rect 251728 378014 252048 378098
rect 251728 377778 251770 378014
rect 252006 377778 252048 378014
rect 251728 377746 252048 377778
rect 246608 374614 246928 374646
rect 246608 374378 246650 374614
rect 246886 374378 246928 374614
rect 246608 374294 246928 374378
rect 246608 374058 246650 374294
rect 246886 374058 246928 374294
rect 246608 374026 246928 374058
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 241488 334894 241808 334926
rect 241488 334658 241530 334894
rect 241766 334658 241808 334894
rect 241488 334574 241808 334658
rect 241488 334338 241530 334574
rect 241766 334338 241808 334574
rect 241488 334306 241808 334338
rect 240114 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 240734 313774
rect 240114 313454 240734 313538
rect 240114 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 240734 313454
rect 236368 295174 236688 295206
rect 236368 294938 236410 295174
rect 236646 294938 236688 295174
rect 236368 294854 236688 294938
rect 236368 294618 236410 294854
rect 236646 294618 236688 294854
rect 236368 294586 236688 294618
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 231248 255454 231568 255486
rect 231248 255218 231290 255454
rect 231526 255218 231568 255454
rect 231248 255134 231568 255218
rect 231248 254898 231290 255134
rect 231526 254898 231568 255134
rect 231248 254866 231568 254898
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 226128 202054 226448 202086
rect 226128 201818 226170 202054
rect 226406 201818 226448 202054
rect 226128 201734 226448 201818
rect 226128 201498 226170 201734
rect 226406 201498 226448 201734
rect 226128 201466 226448 201498
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 228954 194614 229574 230058
rect 232674 234334 233294 269778
rect 240114 277774 240734 313218
rect 243834 317494 244454 352938
rect 253794 363454 254414 398898
rect 257514 403174 258134 438618
rect 264954 446614 265574 482058
rect 268674 486334 269294 521778
rect 276114 529774 276734 565218
rect 279834 569494 280454 604938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 287568 598054 287888 598086
rect 287568 597818 287610 598054
rect 287846 597818 287888 598054
rect 287568 597734 287888 597818
rect 287568 597498 287610 597734
rect 287846 597498 287888 597734
rect 287568 597466 287888 597498
rect 282448 594334 282768 594366
rect 282448 594098 282490 594334
rect 282726 594098 282768 594334
rect 282448 594014 282768 594098
rect 282448 593778 282490 594014
rect 282726 593778 282768 594014
rect 282448 593746 282768 593778
rect 279834 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 280454 569494
rect 279834 569174 280454 569258
rect 279834 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 280454 569174
rect 277328 554614 277648 554646
rect 277328 554378 277370 554614
rect 277606 554378 277648 554614
rect 277328 554294 277648 554378
rect 277328 554058 277370 554294
rect 277606 554058 277648 554294
rect 277328 554026 277648 554058
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 272208 514894 272528 514926
rect 272208 514658 272250 514894
rect 272486 514658 272528 514894
rect 272208 514574 272528 514658
rect 272208 514338 272250 514574
rect 272486 514338 272528 514574
rect 272208 514306 272528 514338
rect 268674 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 269294 486334
rect 268674 486014 269294 486098
rect 268674 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 269294 486014
rect 267088 475174 267408 475206
rect 267088 474938 267130 475174
rect 267366 474938 267408 475174
rect 267088 474854 267408 474938
rect 267088 474618 267130 474854
rect 267366 474618 267408 474854
rect 267088 474586 267408 474618
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 261968 435454 262288 435486
rect 261968 435218 262010 435454
rect 262246 435218 262288 435454
rect 261968 435134 262288 435218
rect 261968 434898 262010 435134
rect 262246 434898 262288 435134
rect 261968 434866 262288 434898
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 256848 382054 257168 382086
rect 256848 381818 256890 382054
rect 257126 381818 257168 382054
rect 256848 381734 257168 381818
rect 256848 381498 256890 381734
rect 257126 381498 257168 381734
rect 256848 381466 257168 381498
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 251728 342334 252048 342366
rect 251728 342098 251770 342334
rect 252006 342098 252048 342334
rect 251728 342014 252048 342098
rect 251728 341778 251770 342014
rect 252006 341778 252048 342014
rect 251728 341746 252048 341778
rect 246608 338614 246928 338646
rect 246608 338378 246650 338614
rect 246886 338378 246928 338614
rect 246608 338294 246928 338378
rect 246608 338058 246650 338294
rect 246886 338058 246928 338294
rect 246608 338026 246928 338058
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 241488 298894 241808 298926
rect 241488 298658 241530 298894
rect 241766 298658 241808 298894
rect 241488 298574 241808 298658
rect 241488 298338 241530 298574
rect 241766 298338 241808 298574
rect 241488 298306 241808 298338
rect 240114 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 240734 277774
rect 240114 277454 240734 277538
rect 240114 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 240734 277454
rect 236368 259174 236688 259206
rect 236368 258938 236410 259174
rect 236646 258938 236688 259174
rect 236368 258854 236688 258938
rect 236368 258618 236410 258854
rect 236646 258618 236688 258854
rect 236368 258586 236688 258618
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 231248 219454 231568 219486
rect 231248 219218 231290 219454
rect 231526 219218 231568 219454
rect 231248 219134 231568 219218
rect 231248 218898 231290 219134
rect 231526 218898 231568 219134
rect 231248 218866 231568 218898
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 226128 166054 226448 166086
rect 226128 165818 226170 166054
rect 226406 165818 226448 166054
rect 226128 165734 226448 165818
rect 226128 165498 226170 165734
rect 226406 165498 226448 165734
rect 226128 165466 226448 165498
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 228954 158614 229574 194058
rect 232674 198334 233294 233778
rect 240114 241774 240734 277218
rect 243834 281494 244454 316938
rect 253794 327454 254414 362898
rect 257514 367174 258134 402618
rect 264954 410614 265574 446058
rect 268674 450334 269294 485778
rect 276114 493774 276734 529218
rect 279834 533494 280454 568938
rect 289794 579454 290414 614898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 602500 297854 622338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 287568 562054 287888 562086
rect 287568 561818 287610 562054
rect 287846 561818 287888 562054
rect 287568 561734 287888 561818
rect 287568 561498 287610 561734
rect 287846 561498 287888 561734
rect 287568 561466 287888 561498
rect 282448 558334 282768 558366
rect 282448 558098 282490 558334
rect 282726 558098 282768 558334
rect 282448 558014 282768 558098
rect 282448 557778 282490 558014
rect 282726 557778 282768 558014
rect 282448 557746 282768 557778
rect 279834 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 280454 533494
rect 279834 533174 280454 533258
rect 279834 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 280454 533174
rect 277328 518614 277648 518646
rect 277328 518378 277370 518614
rect 277606 518378 277648 518614
rect 277328 518294 277648 518378
rect 277328 518058 277370 518294
rect 277606 518058 277648 518294
rect 277328 518026 277648 518058
rect 276114 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 276734 493774
rect 276114 493454 276734 493538
rect 276114 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 276734 493454
rect 272208 478894 272528 478926
rect 272208 478658 272250 478894
rect 272486 478658 272528 478894
rect 272208 478574 272528 478658
rect 272208 478338 272250 478574
rect 272486 478338 272528 478574
rect 272208 478306 272528 478338
rect 268674 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 269294 450334
rect 268674 450014 269294 450098
rect 268674 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 269294 450014
rect 267088 439174 267408 439206
rect 267088 438938 267130 439174
rect 267366 438938 267408 439174
rect 267088 438854 267408 438938
rect 267088 438618 267130 438854
rect 267366 438618 267408 438854
rect 267088 438586 267408 438618
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 261968 399454 262288 399486
rect 261968 399218 262010 399454
rect 262246 399218 262288 399454
rect 261968 399134 262288 399218
rect 261968 398898 262010 399134
rect 262246 398898 262288 399134
rect 261968 398866 262288 398898
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 256848 346054 257168 346086
rect 256848 345818 256890 346054
rect 257126 345818 257168 346054
rect 256848 345734 257168 345818
rect 256848 345498 256890 345734
rect 257126 345498 257168 345734
rect 256848 345466 257168 345498
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 251728 306334 252048 306366
rect 251728 306098 251770 306334
rect 252006 306098 252048 306334
rect 251728 306014 252048 306098
rect 251728 305778 251770 306014
rect 252006 305778 252048 306014
rect 251728 305746 252048 305778
rect 246608 302614 246928 302646
rect 246608 302378 246650 302614
rect 246886 302378 246928 302614
rect 246608 302294 246928 302378
rect 246608 302058 246650 302294
rect 246886 302058 246928 302294
rect 246608 302026 246928 302058
rect 243834 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 244454 281494
rect 243834 281174 244454 281258
rect 243834 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 244454 281174
rect 241488 262894 241808 262926
rect 241488 262658 241530 262894
rect 241766 262658 241808 262894
rect 241488 262574 241808 262658
rect 241488 262338 241530 262574
rect 241766 262338 241808 262574
rect 241488 262306 241808 262338
rect 240114 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 240734 241774
rect 240114 241454 240734 241538
rect 240114 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 240734 241454
rect 236368 223174 236688 223206
rect 236368 222938 236410 223174
rect 236646 222938 236688 223174
rect 236368 222854 236688 222938
rect 236368 222618 236410 222854
rect 236646 222618 236688 222854
rect 236368 222586 236688 222618
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 231248 183454 231568 183486
rect 231248 183218 231290 183454
rect 231526 183218 231568 183454
rect 231248 183134 231568 183218
rect 231248 182898 231290 183134
rect 231526 182898 231568 183134
rect 231248 182866 231568 182898
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 226128 130054 226448 130086
rect 226128 129818 226170 130054
rect 226406 129818 226448 130054
rect 226128 129734 226448 129818
rect 226128 129498 226170 129734
rect 226406 129498 226448 129734
rect 226128 129466 226448 129498
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 228954 122614 229574 158058
rect 232674 162334 233294 197778
rect 240114 205774 240734 241218
rect 243834 245494 244454 280938
rect 253794 291454 254414 326898
rect 257514 331174 258134 366618
rect 264954 374614 265574 410058
rect 268674 414334 269294 449778
rect 276114 457774 276734 493218
rect 279834 497494 280454 532938
rect 289794 543454 290414 578898
rect 292688 579454 293008 579486
rect 292688 579218 292730 579454
rect 292966 579218 293008 579454
rect 292688 579134 293008 579218
rect 292688 578898 292730 579134
rect 292966 578898 293008 579134
rect 292688 578866 293008 578898
rect 293514 547174 294134 582618
rect 297808 583174 298128 583206
rect 297808 582938 297850 583174
rect 298086 582938 298128 583174
rect 297808 582854 298128 582938
rect 297808 582618 297850 582854
rect 298086 582618 298128 582854
rect 297808 582586 298128 582618
rect 300954 554614 301574 590058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 630334 305294 665778
rect 304674 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 305294 630334
rect 304674 630014 305294 630098
rect 304674 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 305294 630014
rect 304674 594334 305294 629778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 602500 309014 633498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 304674 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 305294 594334
rect 304674 594014 305294 594098
rect 304674 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 305294 594014
rect 302928 586894 303248 586926
rect 302928 586658 302970 586894
rect 303206 586658 303248 586894
rect 302928 586574 303248 586658
rect 302928 586338 302970 586574
rect 303206 586338 303248 586574
rect 302928 586306 303248 586338
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 287568 526054 287888 526086
rect 287568 525818 287610 526054
rect 287846 525818 287888 526054
rect 287568 525734 287888 525818
rect 287568 525498 287610 525734
rect 287846 525498 287888 525734
rect 287568 525466 287888 525498
rect 282448 522334 282768 522366
rect 282448 522098 282490 522334
rect 282726 522098 282768 522334
rect 282448 522014 282768 522098
rect 282448 521778 282490 522014
rect 282726 521778 282768 522014
rect 282448 521746 282768 521778
rect 279834 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 280454 497494
rect 279834 497174 280454 497258
rect 279834 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 280454 497174
rect 277328 482614 277648 482646
rect 277328 482378 277370 482614
rect 277606 482378 277648 482614
rect 277328 482294 277648 482378
rect 277328 482058 277370 482294
rect 277606 482058 277648 482294
rect 277328 482026 277648 482058
rect 276114 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 276734 457774
rect 276114 457454 276734 457538
rect 276114 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 276734 457454
rect 272208 442894 272528 442926
rect 272208 442658 272250 442894
rect 272486 442658 272528 442894
rect 272208 442574 272528 442658
rect 272208 442338 272250 442574
rect 272486 442338 272528 442574
rect 272208 442306 272528 442338
rect 268674 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 269294 414334
rect 268674 414014 269294 414098
rect 268674 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 269294 414014
rect 267088 403174 267408 403206
rect 267088 402938 267130 403174
rect 267366 402938 267408 403174
rect 267088 402854 267408 402938
rect 267088 402618 267130 402854
rect 267366 402618 267408 402854
rect 267088 402586 267408 402618
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 261968 363454 262288 363486
rect 261968 363218 262010 363454
rect 262246 363218 262288 363454
rect 261968 363134 262288 363218
rect 261968 362898 262010 363134
rect 262246 362898 262288 363134
rect 261968 362866 262288 362898
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 256848 310054 257168 310086
rect 256848 309818 256890 310054
rect 257126 309818 257168 310054
rect 256848 309734 257168 309818
rect 256848 309498 256890 309734
rect 257126 309498 257168 309734
rect 256848 309466 257168 309498
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 251728 270334 252048 270366
rect 251728 270098 251770 270334
rect 252006 270098 252048 270334
rect 251728 270014 252048 270098
rect 251728 269778 251770 270014
rect 252006 269778 252048 270014
rect 251728 269746 252048 269778
rect 246608 266614 246928 266646
rect 246608 266378 246650 266614
rect 246886 266378 246928 266614
rect 246608 266294 246928 266378
rect 246608 266058 246650 266294
rect 246886 266058 246928 266294
rect 246608 266026 246928 266058
rect 243834 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 244454 245494
rect 243834 245174 244454 245258
rect 243834 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 244454 245174
rect 241488 226894 241808 226926
rect 241488 226658 241530 226894
rect 241766 226658 241808 226894
rect 241488 226574 241808 226658
rect 241488 226338 241530 226574
rect 241766 226338 241808 226574
rect 241488 226306 241808 226338
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 236368 187174 236688 187206
rect 236368 186938 236410 187174
rect 236646 186938 236688 187174
rect 236368 186854 236688 186938
rect 236368 186618 236410 186854
rect 236646 186618 236688 186854
rect 236368 186586 236688 186618
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 231248 147454 231568 147486
rect 231248 147218 231290 147454
rect 231526 147218 231568 147454
rect 231248 147134 231568 147218
rect 231248 146898 231290 147134
rect 231526 146898 231568 147134
rect 231248 146866 231568 146898
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 226128 94054 226448 94086
rect 226128 93818 226170 94054
rect 226406 93818 226448 94054
rect 226128 93734 226448 93818
rect 226128 93498 226170 93734
rect 226406 93498 226448 93734
rect 226128 93466 226448 93498
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 228954 86614 229574 122058
rect 232674 126334 233294 161778
rect 240114 169774 240734 205218
rect 243834 209494 244454 244938
rect 253794 255454 254414 290898
rect 257514 295174 258134 330618
rect 264954 338614 265574 374058
rect 268674 378334 269294 413778
rect 276114 421774 276734 457218
rect 279834 461494 280454 496938
rect 289794 507454 290414 542898
rect 292688 543454 293008 543486
rect 292688 543218 292730 543454
rect 292966 543218 293008 543454
rect 292688 543134 293008 543218
rect 292688 542898 292730 543134
rect 292966 542898 293008 543134
rect 292688 542866 293008 542898
rect 293514 511174 294134 546618
rect 297808 547174 298128 547206
rect 297808 546938 297850 547174
rect 298086 546938 298128 547174
rect 297808 546854 298128 546938
rect 297808 546618 297850 546854
rect 298086 546618 298128 546854
rect 297808 546586 298128 546618
rect 300954 518614 301574 554058
rect 304674 558334 305294 593778
rect 312114 601774 312734 637218
rect 312114 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 312734 601774
rect 312114 601454 312734 601538
rect 312114 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 312734 601454
rect 308048 590614 308368 590646
rect 308048 590378 308090 590614
rect 308326 590378 308368 590614
rect 308048 590294 308368 590378
rect 308048 590058 308090 590294
rect 308326 590058 308368 590294
rect 308048 590026 308368 590058
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 302928 550894 303248 550926
rect 302928 550658 302970 550894
rect 303206 550658 303248 550894
rect 302928 550574 303248 550658
rect 302928 550338 302970 550574
rect 303206 550338 303248 550574
rect 302928 550306 303248 550338
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 287568 490054 287888 490086
rect 287568 489818 287610 490054
rect 287846 489818 287888 490054
rect 287568 489734 287888 489818
rect 287568 489498 287610 489734
rect 287846 489498 287888 489734
rect 287568 489466 287888 489498
rect 282448 486334 282768 486366
rect 282448 486098 282490 486334
rect 282726 486098 282768 486334
rect 282448 486014 282768 486098
rect 282448 485778 282490 486014
rect 282726 485778 282768 486014
rect 282448 485746 282768 485778
rect 279834 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 280454 461494
rect 279834 461174 280454 461258
rect 279834 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 280454 461174
rect 277328 446614 277648 446646
rect 277328 446378 277370 446614
rect 277606 446378 277648 446614
rect 277328 446294 277648 446378
rect 277328 446058 277370 446294
rect 277606 446058 277648 446294
rect 277328 446026 277648 446058
rect 276114 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 276734 421774
rect 276114 421454 276734 421538
rect 276114 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 276734 421454
rect 272208 406894 272528 406926
rect 272208 406658 272250 406894
rect 272486 406658 272528 406894
rect 272208 406574 272528 406658
rect 272208 406338 272250 406574
rect 272486 406338 272528 406574
rect 272208 406306 272528 406338
rect 268674 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 269294 378334
rect 268674 378014 269294 378098
rect 268674 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 269294 378014
rect 267088 367174 267408 367206
rect 267088 366938 267130 367174
rect 267366 366938 267408 367174
rect 267088 366854 267408 366938
rect 267088 366618 267130 366854
rect 267366 366618 267408 366854
rect 267088 366586 267408 366618
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 261968 327454 262288 327486
rect 261968 327218 262010 327454
rect 262246 327218 262288 327454
rect 261968 327134 262288 327218
rect 261968 326898 262010 327134
rect 262246 326898 262288 327134
rect 261968 326866 262288 326898
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 256848 274054 257168 274086
rect 256848 273818 256890 274054
rect 257126 273818 257168 274054
rect 256848 273734 257168 273818
rect 256848 273498 256890 273734
rect 257126 273498 257168 273734
rect 256848 273466 257168 273498
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 251728 234334 252048 234366
rect 251728 234098 251770 234334
rect 252006 234098 252048 234334
rect 251728 234014 252048 234098
rect 251728 233778 251770 234014
rect 252006 233778 252048 234014
rect 251728 233746 252048 233778
rect 246608 230614 246928 230646
rect 246608 230378 246650 230614
rect 246886 230378 246928 230614
rect 246608 230294 246928 230378
rect 246608 230058 246650 230294
rect 246886 230058 246928 230294
rect 246608 230026 246928 230058
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 241488 190894 241808 190926
rect 241488 190658 241530 190894
rect 241766 190658 241808 190894
rect 241488 190574 241808 190658
rect 241488 190338 241530 190574
rect 241766 190338 241808 190574
rect 241488 190306 241808 190338
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 236368 151174 236688 151206
rect 236368 150938 236410 151174
rect 236646 150938 236688 151174
rect 236368 150854 236688 150938
rect 236368 150618 236410 150854
rect 236646 150618 236688 150854
rect 236368 150586 236688 150618
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 231248 111454 231568 111486
rect 231248 111218 231290 111454
rect 231526 111218 231568 111454
rect 231248 111134 231568 111218
rect 231248 110898 231290 111134
rect 231526 110898 231568 111134
rect 231248 110866 231568 110898
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226128 58054 226448 58086
rect 226128 57818 226170 58054
rect 226406 57818 226448 58054
rect 226128 57734 226448 57818
rect 226128 57498 226170 57734
rect 226406 57498 226448 57734
rect 226128 57466 226448 57498
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 228954 50614 229574 86058
rect 232674 90334 233294 125778
rect 240114 133774 240734 169218
rect 243834 173494 244454 208938
rect 253794 219454 254414 254898
rect 257514 259174 258134 294618
rect 264954 302614 265574 338058
rect 268674 342334 269294 377778
rect 276114 385774 276734 421218
rect 279834 425494 280454 460938
rect 289794 471454 290414 506898
rect 292688 507454 293008 507486
rect 292688 507218 292730 507454
rect 292966 507218 293008 507454
rect 292688 507134 293008 507218
rect 292688 506898 292730 507134
rect 292966 506898 293008 507134
rect 292688 506866 293008 506898
rect 293514 475174 294134 510618
rect 297808 511174 298128 511206
rect 297808 510938 297850 511174
rect 298086 510938 298128 511174
rect 297808 510854 298128 510938
rect 297808 510618 297850 510854
rect 298086 510618 298128 510854
rect 297808 510586 298128 510618
rect 300954 482614 301574 518058
rect 304674 522334 305294 557778
rect 312114 565774 312734 601218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 605494 316454 640938
rect 315834 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 316454 605494
rect 315834 605174 316454 605258
rect 315834 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 316454 605174
rect 313168 594334 313488 594366
rect 313168 594098 313210 594334
rect 313446 594098 313488 594334
rect 313168 594014 313488 594098
rect 313168 593778 313210 594014
rect 313446 593778 313488 594014
rect 313168 593746 313488 593778
rect 312114 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 312734 565774
rect 312114 565454 312734 565538
rect 312114 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 312734 565454
rect 308048 554614 308368 554646
rect 308048 554378 308090 554614
rect 308326 554378 308368 554614
rect 308048 554294 308368 554378
rect 308048 554058 308090 554294
rect 308326 554058 308368 554294
rect 308048 554026 308368 554058
rect 304674 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 305294 522334
rect 304674 522014 305294 522098
rect 304674 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 305294 522014
rect 302928 514894 303248 514926
rect 302928 514658 302970 514894
rect 303206 514658 303248 514894
rect 302928 514574 303248 514658
rect 302928 514338 302970 514574
rect 303206 514338 303248 514574
rect 302928 514306 303248 514338
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 287568 454054 287888 454086
rect 287568 453818 287610 454054
rect 287846 453818 287888 454054
rect 287568 453734 287888 453818
rect 287568 453498 287610 453734
rect 287846 453498 287888 453734
rect 287568 453466 287888 453498
rect 282448 450334 282768 450366
rect 282448 450098 282490 450334
rect 282726 450098 282768 450334
rect 282448 450014 282768 450098
rect 282448 449778 282490 450014
rect 282726 449778 282768 450014
rect 282448 449746 282768 449778
rect 279834 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 280454 425494
rect 279834 425174 280454 425258
rect 279834 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 280454 425174
rect 277328 410614 277648 410646
rect 277328 410378 277370 410614
rect 277606 410378 277648 410614
rect 277328 410294 277648 410378
rect 277328 410058 277370 410294
rect 277606 410058 277648 410294
rect 277328 410026 277648 410058
rect 276114 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 276734 385774
rect 276114 385454 276734 385538
rect 276114 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 276734 385454
rect 272208 370894 272528 370926
rect 272208 370658 272250 370894
rect 272486 370658 272528 370894
rect 272208 370574 272528 370658
rect 272208 370338 272250 370574
rect 272486 370338 272528 370574
rect 272208 370306 272528 370338
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 267088 331174 267408 331206
rect 267088 330938 267130 331174
rect 267366 330938 267408 331174
rect 267088 330854 267408 330938
rect 267088 330618 267130 330854
rect 267366 330618 267408 330854
rect 267088 330586 267408 330618
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 261968 291454 262288 291486
rect 261968 291218 262010 291454
rect 262246 291218 262288 291454
rect 261968 291134 262288 291218
rect 261968 290898 262010 291134
rect 262246 290898 262288 291134
rect 261968 290866 262288 290898
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 256848 238054 257168 238086
rect 256848 237818 256890 238054
rect 257126 237818 257168 238054
rect 256848 237734 257168 237818
rect 256848 237498 256890 237734
rect 257126 237498 257168 237734
rect 256848 237466 257168 237498
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 251728 198334 252048 198366
rect 251728 198098 251770 198334
rect 252006 198098 252048 198334
rect 251728 198014 252048 198098
rect 251728 197778 251770 198014
rect 252006 197778 252048 198014
rect 251728 197746 252048 197778
rect 246608 194614 246928 194646
rect 246608 194378 246650 194614
rect 246886 194378 246928 194614
rect 246608 194294 246928 194378
rect 246608 194058 246650 194294
rect 246886 194058 246928 194294
rect 246608 194026 246928 194058
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 241488 154894 241808 154926
rect 241488 154658 241530 154894
rect 241766 154658 241808 154894
rect 241488 154574 241808 154658
rect 241488 154338 241530 154574
rect 241766 154338 241808 154574
rect 241488 154306 241808 154338
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 236368 115174 236688 115206
rect 236368 114938 236410 115174
rect 236646 114938 236688 115174
rect 236368 114854 236688 114938
rect 236368 114618 236410 114854
rect 236646 114618 236688 114854
rect 236368 114586 236688 114618
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 231248 75454 231568 75486
rect 231248 75218 231290 75454
rect 231526 75218 231568 75454
rect 231248 75134 231568 75218
rect 231248 74898 231290 75134
rect 231526 74898 231568 75134
rect 231248 74866 231568 74898
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 226128 22054 226448 22086
rect 226128 21818 226170 22054
rect 226406 21818 226448 22054
rect 226128 21734 226448 21818
rect 226128 21498 226170 21734
rect 226406 21498 226448 21734
rect 226128 21466 226448 21498
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 50058
rect 232674 54334 233294 89778
rect 240114 97774 240734 133218
rect 243834 137494 244454 172938
rect 253794 183454 254414 218898
rect 257514 223174 258134 258618
rect 264954 266614 265574 302058
rect 268674 306334 269294 341778
rect 276114 349774 276734 385218
rect 279834 389494 280454 424938
rect 289794 435454 290414 470898
rect 292688 471454 293008 471486
rect 292688 471218 292730 471454
rect 292966 471218 293008 471454
rect 292688 471134 293008 471218
rect 292688 470898 292730 471134
rect 292966 470898 293008 471134
rect 292688 470866 293008 470898
rect 293514 439174 294134 474618
rect 297808 475174 298128 475206
rect 297808 474938 297850 475174
rect 298086 474938 298128 475174
rect 297808 474854 298128 474938
rect 297808 474618 297850 474854
rect 298086 474618 298128 474854
rect 297808 474586 298128 474618
rect 300954 446614 301574 482058
rect 304674 486334 305294 521778
rect 312114 529774 312734 565218
rect 315834 569494 316454 604938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 318288 598054 318608 598086
rect 318288 597818 318330 598054
rect 318566 597818 318608 598054
rect 318288 597734 318608 597818
rect 318288 597498 318330 597734
rect 318566 597498 318608 597734
rect 318288 597466 318608 597498
rect 323408 579454 323728 579486
rect 323408 579218 323450 579454
rect 323686 579218 323728 579454
rect 323408 579134 323728 579218
rect 323408 578898 323450 579134
rect 323686 578898 323728 579134
rect 323408 578866 323728 578898
rect 325794 579454 326414 614898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 584873 330134 618618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 602500 333854 622338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 630334 341294 665778
rect 340674 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 341294 630334
rect 340674 630014 341294 630098
rect 340674 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 341294 630014
rect 340674 594334 341294 629778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 598054 345014 633498
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 340674 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 341294 594334
rect 340674 594014 341294 594098
rect 340674 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 341294 594014
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 333648 586894 333968 586926
rect 333648 586658 333690 586894
rect 333926 586658 333968 586894
rect 333648 586574 333968 586658
rect 333648 586338 333690 586574
rect 333926 586338 333968 586574
rect 333648 586306 333968 586338
rect 336954 584873 337574 590058
rect 338768 590614 339088 590646
rect 338768 590378 338810 590614
rect 339046 590378 339088 590614
rect 338768 590294 339088 590378
rect 338768 590058 338810 590294
rect 339046 590058 339088 590294
rect 338768 590026 339088 590058
rect 340674 584873 341294 593778
rect 343888 594334 344208 594366
rect 343888 594098 343930 594334
rect 344166 594098 344208 594334
rect 343888 594014 344208 594098
rect 343888 593778 343930 594014
rect 344166 593778 344208 594014
rect 343888 593746 344208 593778
rect 344394 584873 345014 597498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 348114 584873 348734 601218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 349008 598054 349328 598086
rect 349008 597818 349050 598054
rect 349286 597818 349328 598054
rect 349008 597734 349328 597818
rect 349008 597498 349050 597734
rect 349286 597498 349328 597734
rect 349008 597466 349328 597498
rect 351834 584873 352454 604938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 584873 362414 614898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 364368 586894 364688 586926
rect 364368 586658 364410 586894
rect 364646 586658 364688 586894
rect 364368 586574 364688 586658
rect 364368 586338 364410 586574
rect 364646 586338 364688 586574
rect 364368 586306 364688 586338
rect 365514 584873 366134 618618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 602500 369854 622338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 369488 590614 369808 590646
rect 369488 590378 369530 590614
rect 369766 590378 369808 590614
rect 369488 590294 369808 590378
rect 369488 590058 369530 590294
rect 369766 590058 369808 590294
rect 369488 590026 369808 590058
rect 372954 590614 373574 626058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 374608 594334 374928 594366
rect 374608 594098 374650 594334
rect 374886 594098 374928 594334
rect 374608 594014 374928 594098
rect 374608 593778 374650 594014
rect 374886 593778 374928 594014
rect 374608 593746 374928 593778
rect 376674 594334 377294 629778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 379728 598054 380048 598086
rect 379728 597818 379770 598054
rect 380006 597818 380048 598054
rect 379728 597734 380048 597818
rect 379728 597498 379770 597734
rect 380006 597498 380048 597734
rect 379728 597466 380048 597498
rect 380394 598054 381014 633498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 602500 384734 637218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 584873 373574 590058
rect 376674 584873 377294 593778
rect 380394 584873 381014 597498
rect 387834 584873 388454 604938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 395088 586894 395408 586926
rect 395088 586658 395130 586894
rect 395366 586658 395408 586894
rect 395088 586574 395408 586658
rect 395088 586338 395130 586574
rect 395366 586338 395408 586574
rect 395088 586306 395408 586338
rect 397794 584873 398414 614898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 400208 590614 400528 590646
rect 400208 590378 400250 590614
rect 400486 590378 400528 590614
rect 400208 590294 400528 590378
rect 400208 590058 400250 590294
rect 400486 590058 400528 590294
rect 400208 590026 400528 590058
rect 401514 584873 402134 618618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 602500 405854 622338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 405328 594334 405648 594366
rect 405328 594098 405370 594334
rect 405606 594098 405648 594334
rect 405328 594014 405648 594098
rect 405328 593778 405370 594014
rect 405606 593778 405648 594014
rect 405328 593746 405648 593778
rect 408954 590614 409574 626058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 410448 598054 410768 598086
rect 410448 597818 410490 598054
rect 410726 597818 410768 598054
rect 410448 597734 410768 597818
rect 410448 597498 410490 597734
rect 410726 597498 410768 597734
rect 410448 597466 410768 597498
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 584873 409574 590058
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 584873 413294 593778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 602500 420734 637218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 584873 417014 597498
rect 328528 583174 328848 583206
rect 328528 582938 328570 583174
rect 328806 582938 328848 583174
rect 328528 582854 328848 582938
rect 328528 582618 328570 582854
rect 328806 582618 328848 582854
rect 328528 582586 328848 582618
rect 359248 583174 359568 583206
rect 359248 582938 359290 583174
rect 359526 582938 359568 583174
rect 359248 582854 359568 582938
rect 359248 582618 359290 582854
rect 359526 582618 359568 582854
rect 359248 582586 359568 582618
rect 389968 583174 390288 583206
rect 389968 582938 390010 583174
rect 390246 582938 390288 583174
rect 389968 582854 390288 582938
rect 389968 582618 390010 582854
rect 390246 582618 390288 582854
rect 389968 582586 390288 582618
rect 420688 583174 421008 583206
rect 420688 582938 420730 583174
rect 420966 582938 421008 583174
rect 420688 582854 421008 582938
rect 420688 582618 420730 582854
rect 420966 582618 421008 582854
rect 420688 582586 421008 582618
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 315834 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 316454 569494
rect 315834 569174 316454 569258
rect 315834 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 316454 569174
rect 313168 558334 313488 558366
rect 313168 558098 313210 558334
rect 313446 558098 313488 558334
rect 313168 558014 313488 558098
rect 313168 557778 313210 558014
rect 313446 557778 313488 558014
rect 313168 557746 313488 557778
rect 312114 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 312734 529774
rect 312114 529454 312734 529538
rect 312114 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 312734 529454
rect 308048 518614 308368 518646
rect 308048 518378 308090 518614
rect 308326 518378 308368 518614
rect 308048 518294 308368 518378
rect 308048 518058 308090 518294
rect 308326 518058 308368 518294
rect 308048 518026 308368 518058
rect 304674 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 305294 486334
rect 304674 486014 305294 486098
rect 304674 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 305294 486014
rect 302928 478894 303248 478926
rect 302928 478658 302970 478894
rect 303206 478658 303248 478894
rect 302928 478574 303248 478658
rect 302928 478338 302970 478574
rect 303206 478338 303248 478574
rect 302928 478306 303248 478338
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 287568 418054 287888 418086
rect 287568 417818 287610 418054
rect 287846 417818 287888 418054
rect 287568 417734 287888 417818
rect 287568 417498 287610 417734
rect 287846 417498 287888 417734
rect 287568 417466 287888 417498
rect 282448 414334 282768 414366
rect 282448 414098 282490 414334
rect 282726 414098 282768 414334
rect 282448 414014 282768 414098
rect 282448 413778 282490 414014
rect 282726 413778 282768 414014
rect 282448 413746 282768 413778
rect 279834 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 280454 389494
rect 279834 389174 280454 389258
rect 279834 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 280454 389174
rect 277328 374614 277648 374646
rect 277328 374378 277370 374614
rect 277606 374378 277648 374614
rect 277328 374294 277648 374378
rect 277328 374058 277370 374294
rect 277606 374058 277648 374294
rect 277328 374026 277648 374058
rect 276114 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 276734 349774
rect 276114 349454 276734 349538
rect 276114 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 276734 349454
rect 272208 334894 272528 334926
rect 272208 334658 272250 334894
rect 272486 334658 272528 334894
rect 272208 334574 272528 334658
rect 272208 334338 272250 334574
rect 272486 334338 272528 334574
rect 272208 334306 272528 334338
rect 268674 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 269294 306334
rect 268674 306014 269294 306098
rect 268674 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 269294 306014
rect 267088 295174 267408 295206
rect 267088 294938 267130 295174
rect 267366 294938 267408 295174
rect 267088 294854 267408 294938
rect 267088 294618 267130 294854
rect 267366 294618 267408 294854
rect 267088 294586 267408 294618
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 261968 255454 262288 255486
rect 261968 255218 262010 255454
rect 262246 255218 262288 255454
rect 261968 255134 262288 255218
rect 261968 254898 262010 255134
rect 262246 254898 262288 255134
rect 261968 254866 262288 254898
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 256848 202054 257168 202086
rect 256848 201818 256890 202054
rect 257126 201818 257168 202054
rect 256848 201734 257168 201818
rect 256848 201498 256890 201734
rect 257126 201498 257168 201734
rect 256848 201466 257168 201498
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 251728 162334 252048 162366
rect 251728 162098 251770 162334
rect 252006 162098 252048 162334
rect 251728 162014 252048 162098
rect 251728 161778 251770 162014
rect 252006 161778 252048 162014
rect 251728 161746 252048 161778
rect 246608 158614 246928 158646
rect 246608 158378 246650 158614
rect 246886 158378 246928 158614
rect 246608 158294 246928 158378
rect 246608 158058 246650 158294
rect 246886 158058 246928 158294
rect 246608 158026 246928 158058
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 241488 118894 241808 118926
rect 241488 118658 241530 118894
rect 241766 118658 241808 118894
rect 241488 118574 241808 118658
rect 241488 118338 241530 118574
rect 241766 118338 241808 118574
rect 241488 118306 241808 118338
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 236368 79174 236688 79206
rect 236368 78938 236410 79174
rect 236646 78938 236688 79174
rect 236368 78854 236688 78938
rect 236368 78618 236410 78854
rect 236646 78618 236688 78854
rect 236368 78586 236688 78618
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 231248 39454 231568 39486
rect 231248 39218 231290 39454
rect 231526 39218 231568 39454
rect 231248 39134 231568 39218
rect 231248 38898 231290 39134
rect 231526 38898 231568 39134
rect 231248 38866 231568 38898
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 53778
rect 240114 61774 240734 97218
rect 243834 101494 244454 136938
rect 253794 147454 254414 182898
rect 257514 187174 258134 222618
rect 264954 230614 265574 266058
rect 268674 270334 269294 305778
rect 276114 313774 276734 349218
rect 279834 353494 280454 388938
rect 289794 399454 290414 434898
rect 292688 435454 293008 435486
rect 292688 435218 292730 435454
rect 292966 435218 293008 435454
rect 292688 435134 293008 435218
rect 292688 434898 292730 435134
rect 292966 434898 293008 435134
rect 292688 434866 293008 434898
rect 293514 403174 294134 438618
rect 297808 439174 298128 439206
rect 297808 438938 297850 439174
rect 298086 438938 298128 439174
rect 297808 438854 298128 438938
rect 297808 438618 297850 438854
rect 298086 438618 298128 438854
rect 297808 438586 298128 438618
rect 300954 410614 301574 446058
rect 304674 450334 305294 485778
rect 312114 493774 312734 529218
rect 315834 533494 316454 568938
rect 318288 562054 318608 562086
rect 318288 561818 318330 562054
rect 318566 561818 318608 562054
rect 318288 561734 318608 561818
rect 318288 561498 318330 561734
rect 318566 561498 318608 561734
rect 318288 561466 318608 561498
rect 323408 543454 323728 543486
rect 323408 543218 323450 543454
rect 323686 543218 323728 543454
rect 323408 543134 323728 543218
rect 323408 542898 323450 543134
rect 323686 542898 323728 543134
rect 323408 542866 323728 542898
rect 325794 543454 326414 578898
rect 354128 579454 354448 579486
rect 354128 579218 354170 579454
rect 354406 579218 354448 579454
rect 354128 579134 354448 579218
rect 354128 578898 354170 579134
rect 354406 578898 354448 579134
rect 354128 578866 354448 578898
rect 384848 579454 385168 579486
rect 384848 579218 384890 579454
rect 385126 579218 385168 579454
rect 384848 579134 385168 579218
rect 384848 578898 384890 579134
rect 385126 578898 385168 579134
rect 384848 578866 385168 578898
rect 415568 579454 415888 579486
rect 415568 579218 415610 579454
rect 415846 579218 415888 579454
rect 415568 579134 415888 579218
rect 415568 578898 415610 579134
rect 415846 578898 415888 579134
rect 415568 578866 415888 578898
rect 423834 569494 424454 604938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 430928 590614 431248 590646
rect 430928 590378 430970 590614
rect 431206 590378 431248 590614
rect 430928 590294 431248 590378
rect 430928 590058 430970 590294
rect 431206 590058 431248 590294
rect 430928 590026 431248 590058
rect 425808 586894 426128 586926
rect 425808 586658 425850 586894
rect 426086 586658 426128 586894
rect 425808 586574 426128 586658
rect 425808 586338 425850 586574
rect 426086 586338 426128 586574
rect 425808 586306 426128 586338
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 349008 562054 349328 562086
rect 349008 561818 349050 562054
rect 349286 561818 349328 562054
rect 349008 561734 349328 561818
rect 349008 561498 349050 561734
rect 349286 561498 349328 561734
rect 349008 561466 349328 561498
rect 379728 562054 380048 562086
rect 379728 561818 379770 562054
rect 380006 561818 380048 562054
rect 379728 561734 380048 561818
rect 379728 561498 379770 561734
rect 380006 561498 380048 561734
rect 379728 561466 380048 561498
rect 410448 562054 410768 562086
rect 410448 561818 410490 562054
rect 410726 561818 410768 562054
rect 410448 561734 410768 561818
rect 410448 561498 410490 561734
rect 410726 561498 410768 561734
rect 410448 561466 410768 561498
rect 343888 558334 344208 558366
rect 343888 558098 343930 558334
rect 344166 558098 344208 558334
rect 343888 558014 344208 558098
rect 343888 557778 343930 558014
rect 344166 557778 344208 558014
rect 343888 557746 344208 557778
rect 374608 558334 374928 558366
rect 374608 558098 374650 558334
rect 374886 558098 374928 558334
rect 374608 558014 374928 558098
rect 374608 557778 374650 558014
rect 374886 557778 374928 558014
rect 374608 557746 374928 557778
rect 405328 558334 405648 558366
rect 405328 558098 405370 558334
rect 405606 558098 405648 558334
rect 405328 558014 405648 558098
rect 405328 557778 405370 558014
rect 405606 557778 405648 558014
rect 405328 557746 405648 557778
rect 338768 554614 339088 554646
rect 338768 554378 338810 554614
rect 339046 554378 339088 554614
rect 338768 554294 339088 554378
rect 338768 554058 338810 554294
rect 339046 554058 339088 554294
rect 338768 554026 339088 554058
rect 369488 554614 369808 554646
rect 369488 554378 369530 554614
rect 369766 554378 369808 554614
rect 369488 554294 369808 554378
rect 369488 554058 369530 554294
rect 369766 554058 369808 554294
rect 369488 554026 369808 554058
rect 400208 554614 400528 554646
rect 400208 554378 400250 554614
rect 400486 554378 400528 554614
rect 400208 554294 400528 554378
rect 400208 554058 400250 554294
rect 400486 554058 400528 554294
rect 400208 554026 400528 554058
rect 333648 550894 333968 550926
rect 333648 550658 333690 550894
rect 333926 550658 333968 550894
rect 333648 550574 333968 550658
rect 333648 550338 333690 550574
rect 333926 550338 333968 550574
rect 333648 550306 333968 550338
rect 364368 550894 364688 550926
rect 364368 550658 364410 550894
rect 364646 550658 364688 550894
rect 364368 550574 364688 550658
rect 364368 550338 364410 550574
rect 364646 550338 364688 550574
rect 364368 550306 364688 550338
rect 395088 550894 395408 550926
rect 395088 550658 395130 550894
rect 395366 550658 395408 550894
rect 395088 550574 395408 550658
rect 395088 550338 395130 550574
rect 395366 550338 395408 550574
rect 395088 550306 395408 550338
rect 328528 547174 328848 547206
rect 328528 546938 328570 547174
rect 328806 546938 328848 547174
rect 328528 546854 328848 546938
rect 328528 546618 328570 546854
rect 328806 546618 328848 546854
rect 328528 546586 328848 546618
rect 359248 547174 359568 547206
rect 359248 546938 359290 547174
rect 359526 546938 359568 547174
rect 359248 546854 359568 546938
rect 359248 546618 359290 546854
rect 359526 546618 359568 546854
rect 359248 546586 359568 546618
rect 389968 547174 390288 547206
rect 389968 546938 390010 547174
rect 390246 546938 390288 547174
rect 389968 546854 390288 546938
rect 389968 546618 390010 546854
rect 390246 546618 390288 546854
rect 389968 546586 390288 546618
rect 420688 547174 421008 547206
rect 420688 546938 420730 547174
rect 420966 546938 421008 547174
rect 420688 546854 421008 546938
rect 420688 546618 420730 546854
rect 420966 546618 421008 546854
rect 420688 546586 421008 546618
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 315834 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 316454 533494
rect 315834 533174 316454 533258
rect 315834 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 316454 533174
rect 313168 522334 313488 522366
rect 313168 522098 313210 522334
rect 313446 522098 313488 522334
rect 313168 522014 313488 522098
rect 313168 521778 313210 522014
rect 313446 521778 313488 522014
rect 313168 521746 313488 521778
rect 312114 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 312734 493774
rect 312114 493454 312734 493538
rect 312114 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 312734 493454
rect 308048 482614 308368 482646
rect 308048 482378 308090 482614
rect 308326 482378 308368 482614
rect 308048 482294 308368 482378
rect 308048 482058 308090 482294
rect 308326 482058 308368 482294
rect 308048 482026 308368 482058
rect 304674 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 305294 450334
rect 304674 450014 305294 450098
rect 304674 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 305294 450014
rect 302928 442894 303248 442926
rect 302928 442658 302970 442894
rect 303206 442658 303248 442894
rect 302928 442574 303248 442658
rect 302928 442338 302970 442574
rect 303206 442338 303248 442574
rect 302928 442306 303248 442338
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 287568 382054 287888 382086
rect 287568 381818 287610 382054
rect 287846 381818 287888 382054
rect 287568 381734 287888 381818
rect 287568 381498 287610 381734
rect 287846 381498 287888 381734
rect 287568 381466 287888 381498
rect 282448 378334 282768 378366
rect 282448 378098 282490 378334
rect 282726 378098 282768 378334
rect 282448 378014 282768 378098
rect 282448 377778 282490 378014
rect 282726 377778 282768 378014
rect 282448 377746 282768 377778
rect 279834 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 280454 353494
rect 279834 353174 280454 353258
rect 279834 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 280454 353174
rect 277328 338614 277648 338646
rect 277328 338378 277370 338614
rect 277606 338378 277648 338614
rect 277328 338294 277648 338378
rect 277328 338058 277370 338294
rect 277606 338058 277648 338294
rect 277328 338026 277648 338058
rect 276114 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 276734 313774
rect 276114 313454 276734 313538
rect 276114 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 276734 313454
rect 272208 298894 272528 298926
rect 272208 298658 272250 298894
rect 272486 298658 272528 298894
rect 272208 298574 272528 298658
rect 272208 298338 272250 298574
rect 272486 298338 272528 298574
rect 272208 298306 272528 298338
rect 268674 270098 268706 270334
rect 268942 270098 269026 270334
rect 269262 270098 269294 270334
rect 268674 270014 269294 270098
rect 268674 269778 268706 270014
rect 268942 269778 269026 270014
rect 269262 269778 269294 270014
rect 267088 259174 267408 259206
rect 267088 258938 267130 259174
rect 267366 258938 267408 259174
rect 267088 258854 267408 258938
rect 267088 258618 267130 258854
rect 267366 258618 267408 258854
rect 267088 258586 267408 258618
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 261968 219454 262288 219486
rect 261968 219218 262010 219454
rect 262246 219218 262288 219454
rect 261968 219134 262288 219218
rect 261968 218898 262010 219134
rect 262246 218898 262288 219134
rect 261968 218866 262288 218898
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 256848 166054 257168 166086
rect 256848 165818 256890 166054
rect 257126 165818 257168 166054
rect 256848 165734 257168 165818
rect 256848 165498 256890 165734
rect 257126 165498 257168 165734
rect 256848 165466 257168 165498
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 251728 126334 252048 126366
rect 251728 126098 251770 126334
rect 252006 126098 252048 126334
rect 251728 126014 252048 126098
rect 251728 125778 251770 126014
rect 252006 125778 252048 126014
rect 251728 125746 252048 125778
rect 246608 122614 246928 122646
rect 246608 122378 246650 122614
rect 246886 122378 246928 122614
rect 246608 122294 246928 122378
rect 246608 122058 246650 122294
rect 246886 122058 246928 122294
rect 246608 122026 246928 122058
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 241488 82894 241808 82926
rect 241488 82658 241530 82894
rect 241766 82658 241808 82894
rect 241488 82574 241808 82658
rect 241488 82338 241530 82574
rect 241766 82338 241808 82574
rect 241488 82306 241808 82338
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 236368 43174 236688 43206
rect 236368 42938 236410 43174
rect 236646 42938 236688 43174
rect 236368 42854 236688 42938
rect 236368 42618 236410 42854
rect 236646 42618 236688 42854
rect 236368 42586 236688 42618
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 240114 25774 240734 61218
rect 243834 65494 244454 100938
rect 253794 111454 254414 146898
rect 257514 151174 258134 186618
rect 264954 194614 265574 230058
rect 268674 234334 269294 269778
rect 276114 277774 276734 313218
rect 279834 317494 280454 352938
rect 289794 363454 290414 398898
rect 292688 399454 293008 399486
rect 292688 399218 292730 399454
rect 292966 399218 293008 399454
rect 292688 399134 293008 399218
rect 292688 398898 292730 399134
rect 292966 398898 293008 399134
rect 292688 398866 293008 398898
rect 293514 367174 294134 402618
rect 297808 403174 298128 403206
rect 297808 402938 297850 403174
rect 298086 402938 298128 403174
rect 297808 402854 298128 402938
rect 297808 402618 297850 402854
rect 298086 402618 298128 402854
rect 297808 402586 298128 402618
rect 300954 374614 301574 410058
rect 304674 414334 305294 449778
rect 312114 457774 312734 493218
rect 315834 497494 316454 532938
rect 318288 526054 318608 526086
rect 318288 525818 318330 526054
rect 318566 525818 318608 526054
rect 318288 525734 318608 525818
rect 318288 525498 318330 525734
rect 318566 525498 318608 525734
rect 318288 525466 318608 525498
rect 323408 507454 323728 507486
rect 323408 507218 323450 507454
rect 323686 507218 323728 507454
rect 323408 507134 323728 507218
rect 323408 506898 323450 507134
rect 323686 506898 323728 507134
rect 323408 506866 323728 506898
rect 325794 507454 326414 542898
rect 354128 543454 354448 543486
rect 354128 543218 354170 543454
rect 354406 543218 354448 543454
rect 354128 543134 354448 543218
rect 354128 542898 354170 543134
rect 354406 542898 354448 543134
rect 354128 542866 354448 542898
rect 384848 543454 385168 543486
rect 384848 543218 384890 543454
rect 385126 543218 385168 543454
rect 384848 543134 385168 543218
rect 384848 542898 384890 543134
rect 385126 542898 385168 543134
rect 384848 542866 385168 542898
rect 415568 543454 415888 543486
rect 415568 543218 415610 543454
rect 415846 543218 415888 543454
rect 415568 543134 415888 543218
rect 415568 542898 415610 543134
rect 415846 542898 415888 543134
rect 415568 542866 415888 542898
rect 423834 533494 424454 568938
rect 433794 579454 434414 614898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 436048 594334 436368 594366
rect 436048 594098 436090 594334
rect 436326 594098 436368 594334
rect 436048 594014 436368 594098
rect 436048 593778 436090 594014
rect 436326 593778 436368 594014
rect 436048 593746 436368 593778
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 430928 554614 431248 554646
rect 430928 554378 430970 554614
rect 431206 554378 431248 554614
rect 430928 554294 431248 554378
rect 430928 554058 430970 554294
rect 431206 554058 431248 554294
rect 430928 554026 431248 554058
rect 425808 550894 426128 550926
rect 425808 550658 425850 550894
rect 426086 550658 426128 550894
rect 425808 550574 426128 550658
rect 425808 550338 425850 550574
rect 426086 550338 426128 550574
rect 425808 550306 426128 550338
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 349008 526054 349328 526086
rect 349008 525818 349050 526054
rect 349286 525818 349328 526054
rect 349008 525734 349328 525818
rect 349008 525498 349050 525734
rect 349286 525498 349328 525734
rect 349008 525466 349328 525498
rect 379728 526054 380048 526086
rect 379728 525818 379770 526054
rect 380006 525818 380048 526054
rect 379728 525734 380048 525818
rect 379728 525498 379770 525734
rect 380006 525498 380048 525734
rect 379728 525466 380048 525498
rect 410448 526054 410768 526086
rect 410448 525818 410490 526054
rect 410726 525818 410768 526054
rect 410448 525734 410768 525818
rect 410448 525498 410490 525734
rect 410726 525498 410768 525734
rect 410448 525466 410768 525498
rect 343888 522334 344208 522366
rect 343888 522098 343930 522334
rect 344166 522098 344208 522334
rect 343888 522014 344208 522098
rect 343888 521778 343930 522014
rect 344166 521778 344208 522014
rect 343888 521746 344208 521778
rect 374608 522334 374928 522366
rect 374608 522098 374650 522334
rect 374886 522098 374928 522334
rect 374608 522014 374928 522098
rect 374608 521778 374650 522014
rect 374886 521778 374928 522014
rect 374608 521746 374928 521778
rect 405328 522334 405648 522366
rect 405328 522098 405370 522334
rect 405606 522098 405648 522334
rect 405328 522014 405648 522098
rect 405328 521778 405370 522014
rect 405606 521778 405648 522014
rect 405328 521746 405648 521778
rect 338768 518614 339088 518646
rect 338768 518378 338810 518614
rect 339046 518378 339088 518614
rect 338768 518294 339088 518378
rect 338768 518058 338810 518294
rect 339046 518058 339088 518294
rect 338768 518026 339088 518058
rect 369488 518614 369808 518646
rect 369488 518378 369530 518614
rect 369766 518378 369808 518614
rect 369488 518294 369808 518378
rect 369488 518058 369530 518294
rect 369766 518058 369808 518294
rect 369488 518026 369808 518058
rect 400208 518614 400528 518646
rect 400208 518378 400250 518614
rect 400486 518378 400528 518614
rect 400208 518294 400528 518378
rect 400208 518058 400250 518294
rect 400486 518058 400528 518294
rect 400208 518026 400528 518058
rect 333648 514894 333968 514926
rect 333648 514658 333690 514894
rect 333926 514658 333968 514894
rect 333648 514574 333968 514658
rect 333648 514338 333690 514574
rect 333926 514338 333968 514574
rect 333648 514306 333968 514338
rect 364368 514894 364688 514926
rect 364368 514658 364410 514894
rect 364646 514658 364688 514894
rect 364368 514574 364688 514658
rect 364368 514338 364410 514574
rect 364646 514338 364688 514574
rect 364368 514306 364688 514338
rect 395088 514894 395408 514926
rect 395088 514658 395130 514894
rect 395366 514658 395408 514894
rect 395088 514574 395408 514658
rect 395088 514338 395130 514574
rect 395366 514338 395408 514574
rect 395088 514306 395408 514338
rect 328528 511174 328848 511206
rect 328528 510938 328570 511174
rect 328806 510938 328848 511174
rect 328528 510854 328848 510938
rect 328528 510618 328570 510854
rect 328806 510618 328848 510854
rect 328528 510586 328848 510618
rect 359248 511174 359568 511206
rect 359248 510938 359290 511174
rect 359526 510938 359568 511174
rect 359248 510854 359568 510938
rect 359248 510618 359290 510854
rect 359526 510618 359568 510854
rect 359248 510586 359568 510618
rect 389968 511174 390288 511206
rect 389968 510938 390010 511174
rect 390246 510938 390288 511174
rect 389968 510854 390288 510938
rect 389968 510618 390010 510854
rect 390246 510618 390288 510854
rect 389968 510586 390288 510618
rect 420688 511174 421008 511206
rect 420688 510938 420730 511174
rect 420966 510938 421008 511174
rect 420688 510854 421008 510938
rect 420688 510618 420730 510854
rect 420966 510618 421008 510854
rect 420688 510586 421008 510618
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 315834 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 316454 497494
rect 315834 497174 316454 497258
rect 315834 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 316454 497174
rect 313168 486334 313488 486366
rect 313168 486098 313210 486334
rect 313446 486098 313488 486334
rect 313168 486014 313488 486098
rect 313168 485778 313210 486014
rect 313446 485778 313488 486014
rect 313168 485746 313488 485778
rect 312114 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 312734 457774
rect 312114 457454 312734 457538
rect 312114 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 312734 457454
rect 308048 446614 308368 446646
rect 308048 446378 308090 446614
rect 308326 446378 308368 446614
rect 308048 446294 308368 446378
rect 308048 446058 308090 446294
rect 308326 446058 308368 446294
rect 308048 446026 308368 446058
rect 304674 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 305294 414334
rect 304674 414014 305294 414098
rect 304674 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 305294 414014
rect 302928 406894 303248 406926
rect 302928 406658 302970 406894
rect 303206 406658 303248 406894
rect 302928 406574 303248 406658
rect 302928 406338 302970 406574
rect 303206 406338 303248 406574
rect 302928 406306 303248 406338
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 287568 346054 287888 346086
rect 287568 345818 287610 346054
rect 287846 345818 287888 346054
rect 287568 345734 287888 345818
rect 287568 345498 287610 345734
rect 287846 345498 287888 345734
rect 287568 345466 287888 345498
rect 282448 342334 282768 342366
rect 282448 342098 282490 342334
rect 282726 342098 282768 342334
rect 282448 342014 282768 342098
rect 282448 341778 282490 342014
rect 282726 341778 282768 342014
rect 282448 341746 282768 341778
rect 279834 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 280454 317494
rect 279834 317174 280454 317258
rect 279834 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 280454 317174
rect 277328 302614 277648 302646
rect 277328 302378 277370 302614
rect 277606 302378 277648 302614
rect 277328 302294 277648 302378
rect 277328 302058 277370 302294
rect 277606 302058 277648 302294
rect 277328 302026 277648 302058
rect 276114 277538 276146 277774
rect 276382 277538 276466 277774
rect 276702 277538 276734 277774
rect 276114 277454 276734 277538
rect 276114 277218 276146 277454
rect 276382 277218 276466 277454
rect 276702 277218 276734 277454
rect 272208 262894 272528 262926
rect 272208 262658 272250 262894
rect 272486 262658 272528 262894
rect 272208 262574 272528 262658
rect 272208 262338 272250 262574
rect 272486 262338 272528 262574
rect 272208 262306 272528 262338
rect 268674 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 269294 234334
rect 268674 234014 269294 234098
rect 268674 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 269294 234014
rect 267088 223174 267408 223206
rect 267088 222938 267130 223174
rect 267366 222938 267408 223174
rect 267088 222854 267408 222938
rect 267088 222618 267130 222854
rect 267366 222618 267408 222854
rect 267088 222586 267408 222618
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 261968 183454 262288 183486
rect 261968 183218 262010 183454
rect 262246 183218 262288 183454
rect 261968 183134 262288 183218
rect 261968 182898 262010 183134
rect 262246 182898 262288 183134
rect 261968 182866 262288 182898
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 256848 130054 257168 130086
rect 256848 129818 256890 130054
rect 257126 129818 257168 130054
rect 256848 129734 257168 129818
rect 256848 129498 256890 129734
rect 257126 129498 257168 129734
rect 256848 129466 257168 129498
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 251728 90334 252048 90366
rect 251728 90098 251770 90334
rect 252006 90098 252048 90334
rect 251728 90014 252048 90098
rect 251728 89778 251770 90014
rect 252006 89778 252048 90014
rect 251728 89746 252048 89778
rect 246608 86614 246928 86646
rect 246608 86378 246650 86614
rect 246886 86378 246928 86614
rect 246608 86294 246928 86378
rect 246608 86058 246650 86294
rect 246886 86058 246928 86294
rect 246608 86026 246928 86058
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 241488 46894 241808 46926
rect 241488 46658 241530 46894
rect 241766 46658 241808 46894
rect 241488 46574 241808 46658
rect 241488 46338 241530 46574
rect 241766 46338 241808 46574
rect 241488 46306 241808 46338
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 236368 7174 236688 7206
rect 236368 6938 236410 7174
rect 236646 6938 236688 7174
rect 236368 6854 236688 6938
rect 236368 6618 236410 6854
rect 236646 6618 236688 6854
rect 236368 6586 236688 6618
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 -5146 237014 2988
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 -6106 240734 25218
rect 243834 29494 244454 64938
rect 253794 75454 254414 110898
rect 257514 115174 258134 150618
rect 264954 158614 265574 194058
rect 268674 198334 269294 233778
rect 276114 241774 276734 277218
rect 279834 281494 280454 316938
rect 289794 327454 290414 362898
rect 292688 363454 293008 363486
rect 292688 363218 292730 363454
rect 292966 363218 293008 363454
rect 292688 363134 293008 363218
rect 292688 362898 292730 363134
rect 292966 362898 293008 363134
rect 292688 362866 293008 362898
rect 293514 331174 294134 366618
rect 297808 367174 298128 367206
rect 297808 366938 297850 367174
rect 298086 366938 298128 367174
rect 297808 366854 298128 366938
rect 297808 366618 297850 366854
rect 298086 366618 298128 366854
rect 297808 366586 298128 366618
rect 300954 338614 301574 374058
rect 304674 378334 305294 413778
rect 312114 421774 312734 457218
rect 315834 461494 316454 496938
rect 318288 490054 318608 490086
rect 318288 489818 318330 490054
rect 318566 489818 318608 490054
rect 318288 489734 318608 489818
rect 318288 489498 318330 489734
rect 318566 489498 318608 489734
rect 318288 489466 318608 489498
rect 323408 471454 323728 471486
rect 323408 471218 323450 471454
rect 323686 471218 323728 471454
rect 323408 471134 323728 471218
rect 323408 470898 323450 471134
rect 323686 470898 323728 471134
rect 323408 470866 323728 470898
rect 325794 471454 326414 506898
rect 354128 507454 354448 507486
rect 354128 507218 354170 507454
rect 354406 507218 354448 507454
rect 354128 507134 354448 507218
rect 354128 506898 354170 507134
rect 354406 506898 354448 507134
rect 354128 506866 354448 506898
rect 384848 507454 385168 507486
rect 384848 507218 384890 507454
rect 385126 507218 385168 507454
rect 384848 507134 385168 507218
rect 384848 506898 384890 507134
rect 385126 506898 385168 507134
rect 384848 506866 385168 506898
rect 415568 507454 415888 507486
rect 415568 507218 415610 507454
rect 415846 507218 415888 507454
rect 415568 507134 415888 507218
rect 415568 506898 415610 507134
rect 415846 506898 415888 507134
rect 415568 506866 415888 506898
rect 423834 497494 424454 532938
rect 433794 543454 434414 578898
rect 437514 583174 438134 618618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 602500 441854 622338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 441168 598054 441488 598086
rect 441168 597818 441210 598054
rect 441446 597818 441488 598054
rect 441168 597734 441488 597818
rect 441168 597498 441210 597734
rect 441446 597498 441488 597734
rect 441168 597466 441488 597498
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 436048 558334 436368 558366
rect 436048 558098 436090 558334
rect 436326 558098 436368 558334
rect 436048 558014 436368 558098
rect 436048 557778 436090 558014
rect 436326 557778 436368 558014
rect 436048 557746 436368 557778
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 430928 518614 431248 518646
rect 430928 518378 430970 518614
rect 431206 518378 431248 518614
rect 430928 518294 431248 518378
rect 430928 518058 430970 518294
rect 431206 518058 431248 518294
rect 430928 518026 431248 518058
rect 425808 514894 426128 514926
rect 425808 514658 425850 514894
rect 426086 514658 426128 514894
rect 425808 514574 426128 514658
rect 425808 514338 425850 514574
rect 426086 514338 426128 514574
rect 425808 514306 426128 514338
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 349008 490054 349328 490086
rect 349008 489818 349050 490054
rect 349286 489818 349328 490054
rect 349008 489734 349328 489818
rect 349008 489498 349050 489734
rect 349286 489498 349328 489734
rect 349008 489466 349328 489498
rect 379728 490054 380048 490086
rect 379728 489818 379770 490054
rect 380006 489818 380048 490054
rect 379728 489734 380048 489818
rect 379728 489498 379770 489734
rect 380006 489498 380048 489734
rect 379728 489466 380048 489498
rect 410448 490054 410768 490086
rect 410448 489818 410490 490054
rect 410726 489818 410768 490054
rect 410448 489734 410768 489818
rect 410448 489498 410490 489734
rect 410726 489498 410768 489734
rect 410448 489466 410768 489498
rect 343888 486334 344208 486366
rect 343888 486098 343930 486334
rect 344166 486098 344208 486334
rect 343888 486014 344208 486098
rect 343888 485778 343930 486014
rect 344166 485778 344208 486014
rect 343888 485746 344208 485778
rect 374608 486334 374928 486366
rect 374608 486098 374650 486334
rect 374886 486098 374928 486334
rect 374608 486014 374928 486098
rect 374608 485778 374650 486014
rect 374886 485778 374928 486014
rect 374608 485746 374928 485778
rect 405328 486334 405648 486366
rect 405328 486098 405370 486334
rect 405606 486098 405648 486334
rect 405328 486014 405648 486098
rect 405328 485778 405370 486014
rect 405606 485778 405648 486014
rect 405328 485746 405648 485778
rect 338768 482614 339088 482646
rect 338768 482378 338810 482614
rect 339046 482378 339088 482614
rect 338768 482294 339088 482378
rect 338768 482058 338810 482294
rect 339046 482058 339088 482294
rect 338768 482026 339088 482058
rect 369488 482614 369808 482646
rect 369488 482378 369530 482614
rect 369766 482378 369808 482614
rect 369488 482294 369808 482378
rect 369488 482058 369530 482294
rect 369766 482058 369808 482294
rect 369488 482026 369808 482058
rect 400208 482614 400528 482646
rect 400208 482378 400250 482614
rect 400486 482378 400528 482614
rect 400208 482294 400528 482378
rect 400208 482058 400250 482294
rect 400486 482058 400528 482294
rect 400208 482026 400528 482058
rect 333648 478894 333968 478926
rect 333648 478658 333690 478894
rect 333926 478658 333968 478894
rect 333648 478574 333968 478658
rect 333648 478338 333690 478574
rect 333926 478338 333968 478574
rect 333648 478306 333968 478338
rect 364368 478894 364688 478926
rect 364368 478658 364410 478894
rect 364646 478658 364688 478894
rect 364368 478574 364688 478658
rect 364368 478338 364410 478574
rect 364646 478338 364688 478574
rect 364368 478306 364688 478338
rect 395088 478894 395408 478926
rect 395088 478658 395130 478894
rect 395366 478658 395408 478894
rect 395088 478574 395408 478658
rect 395088 478338 395130 478574
rect 395366 478338 395408 478574
rect 395088 478306 395408 478338
rect 328528 475174 328848 475206
rect 328528 474938 328570 475174
rect 328806 474938 328848 475174
rect 328528 474854 328848 474938
rect 328528 474618 328570 474854
rect 328806 474618 328848 474854
rect 328528 474586 328848 474618
rect 359248 475174 359568 475206
rect 359248 474938 359290 475174
rect 359526 474938 359568 475174
rect 359248 474854 359568 474938
rect 359248 474618 359290 474854
rect 359526 474618 359568 474854
rect 359248 474586 359568 474618
rect 389968 475174 390288 475206
rect 389968 474938 390010 475174
rect 390246 474938 390288 475174
rect 389968 474854 390288 474938
rect 389968 474618 390010 474854
rect 390246 474618 390288 474854
rect 389968 474586 390288 474618
rect 420688 475174 421008 475206
rect 420688 474938 420730 475174
rect 420966 474938 421008 475174
rect 420688 474854 421008 474938
rect 420688 474618 420730 474854
rect 420966 474618 421008 474854
rect 420688 474586 421008 474618
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 315834 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 316454 461494
rect 315834 461174 316454 461258
rect 315834 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 316454 461174
rect 313168 450334 313488 450366
rect 313168 450098 313210 450334
rect 313446 450098 313488 450334
rect 313168 450014 313488 450098
rect 313168 449778 313210 450014
rect 313446 449778 313488 450014
rect 313168 449746 313488 449778
rect 312114 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 312734 421774
rect 312114 421454 312734 421538
rect 312114 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 312734 421454
rect 308048 410614 308368 410646
rect 308048 410378 308090 410614
rect 308326 410378 308368 410614
rect 308048 410294 308368 410378
rect 308048 410058 308090 410294
rect 308326 410058 308368 410294
rect 308048 410026 308368 410058
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 302928 370894 303248 370926
rect 302928 370658 302970 370894
rect 303206 370658 303248 370894
rect 302928 370574 303248 370658
rect 302928 370338 302970 370574
rect 303206 370338 303248 370574
rect 302928 370306 303248 370338
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 287568 310054 287888 310086
rect 287568 309818 287610 310054
rect 287846 309818 287888 310054
rect 287568 309734 287888 309818
rect 287568 309498 287610 309734
rect 287846 309498 287888 309734
rect 287568 309466 287888 309498
rect 282448 306334 282768 306366
rect 282448 306098 282490 306334
rect 282726 306098 282768 306334
rect 282448 306014 282768 306098
rect 282448 305778 282490 306014
rect 282726 305778 282768 306014
rect 282448 305746 282768 305778
rect 279834 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 280454 281494
rect 279834 281174 280454 281258
rect 279834 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 280454 281174
rect 277328 266614 277648 266646
rect 277328 266378 277370 266614
rect 277606 266378 277648 266614
rect 277328 266294 277648 266378
rect 277328 266058 277370 266294
rect 277606 266058 277648 266294
rect 277328 266026 277648 266058
rect 276114 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 276734 241774
rect 276114 241454 276734 241538
rect 276114 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 276734 241454
rect 272208 226894 272528 226926
rect 272208 226658 272250 226894
rect 272486 226658 272528 226894
rect 272208 226574 272528 226658
rect 272208 226338 272250 226574
rect 272486 226338 272528 226574
rect 272208 226306 272528 226338
rect 268674 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 269294 198334
rect 268674 198014 269294 198098
rect 268674 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 269294 198014
rect 267088 187174 267408 187206
rect 267088 186938 267130 187174
rect 267366 186938 267408 187174
rect 267088 186854 267408 186938
rect 267088 186618 267130 186854
rect 267366 186618 267408 186854
rect 267088 186586 267408 186618
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 261968 147454 262288 147486
rect 261968 147218 262010 147454
rect 262246 147218 262288 147454
rect 261968 147134 262288 147218
rect 261968 146898 262010 147134
rect 262246 146898 262288 147134
rect 261968 146866 262288 146898
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 256848 94054 257168 94086
rect 256848 93818 256890 94054
rect 257126 93818 257168 94054
rect 256848 93734 257168 93818
rect 256848 93498 256890 93734
rect 257126 93498 257168 93734
rect 256848 93466 257168 93498
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 251728 54334 252048 54366
rect 251728 54098 251770 54334
rect 252006 54098 252048 54334
rect 251728 54014 252048 54098
rect 251728 53778 251770 54014
rect 252006 53778 252048 54014
rect 251728 53746 252048 53778
rect 246608 50614 246928 50646
rect 246608 50378 246650 50614
rect 246886 50378 246928 50614
rect 246608 50294 246928 50378
rect 246608 50058 246650 50294
rect 246886 50058 246928 50294
rect 246608 50026 246928 50058
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 241488 10894 241808 10926
rect 241488 10658 241530 10894
rect 241766 10658 241808 10894
rect 241488 10574 241808 10658
rect 241488 10338 241530 10574
rect 241766 10338 241808 10574
rect 241488 10306 241808 10338
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 -7066 244454 28938
rect 253794 39454 254414 74898
rect 257514 79174 258134 114618
rect 264954 122614 265574 158058
rect 268674 162334 269294 197778
rect 276114 205774 276734 241218
rect 279834 245494 280454 280938
rect 289794 291454 290414 326898
rect 292688 327454 293008 327486
rect 292688 327218 292730 327454
rect 292966 327218 293008 327454
rect 292688 327134 293008 327218
rect 292688 326898 292730 327134
rect 292966 326898 293008 327134
rect 292688 326866 293008 326898
rect 293514 295174 294134 330618
rect 297808 331174 298128 331206
rect 297808 330938 297850 331174
rect 298086 330938 298128 331174
rect 297808 330854 298128 330938
rect 297808 330618 297850 330854
rect 298086 330618 298128 330854
rect 297808 330586 298128 330618
rect 300954 302614 301574 338058
rect 304674 342334 305294 377778
rect 312114 385774 312734 421218
rect 315834 425494 316454 460938
rect 318288 454054 318608 454086
rect 318288 453818 318330 454054
rect 318566 453818 318608 454054
rect 318288 453734 318608 453818
rect 318288 453498 318330 453734
rect 318566 453498 318608 453734
rect 318288 453466 318608 453498
rect 323408 435454 323728 435486
rect 323408 435218 323450 435454
rect 323686 435218 323728 435454
rect 323408 435134 323728 435218
rect 323408 434898 323450 435134
rect 323686 434898 323728 435134
rect 323408 434866 323728 434898
rect 325794 435454 326414 470898
rect 354128 471454 354448 471486
rect 354128 471218 354170 471454
rect 354406 471218 354448 471454
rect 354128 471134 354448 471218
rect 354128 470898 354170 471134
rect 354406 470898 354448 471134
rect 354128 470866 354448 470898
rect 384848 471454 385168 471486
rect 384848 471218 384890 471454
rect 385126 471218 385168 471454
rect 384848 471134 385168 471218
rect 384848 470898 384890 471134
rect 385126 470898 385168 471134
rect 384848 470866 385168 470898
rect 415568 471454 415888 471486
rect 415568 471218 415610 471454
rect 415846 471218 415888 471454
rect 415568 471134 415888 471218
rect 415568 470898 415610 471134
rect 415846 470898 415888 471134
rect 415568 470866 415888 470898
rect 423834 461494 424454 496938
rect 433794 507454 434414 542898
rect 437514 547174 438134 582618
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 441168 562054 441488 562086
rect 441168 561818 441210 562054
rect 441446 561818 441488 562054
rect 441168 561734 441488 561818
rect 441168 561498 441210 561734
rect 441446 561498 441488 561734
rect 441168 561466 441488 561498
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 436048 522334 436368 522366
rect 436048 522098 436090 522334
rect 436326 522098 436368 522334
rect 436048 522014 436368 522098
rect 436048 521778 436090 522014
rect 436326 521778 436368 522014
rect 436048 521746 436368 521778
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 430928 482614 431248 482646
rect 430928 482378 430970 482614
rect 431206 482378 431248 482614
rect 430928 482294 431248 482378
rect 430928 482058 430970 482294
rect 431206 482058 431248 482294
rect 430928 482026 431248 482058
rect 425808 478894 426128 478926
rect 425808 478658 425850 478894
rect 426086 478658 426128 478894
rect 425808 478574 426128 478658
rect 425808 478338 425850 478574
rect 426086 478338 426128 478574
rect 425808 478306 426128 478338
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 349008 454054 349328 454086
rect 349008 453818 349050 454054
rect 349286 453818 349328 454054
rect 349008 453734 349328 453818
rect 349008 453498 349050 453734
rect 349286 453498 349328 453734
rect 349008 453466 349328 453498
rect 379728 454054 380048 454086
rect 379728 453818 379770 454054
rect 380006 453818 380048 454054
rect 379728 453734 380048 453818
rect 379728 453498 379770 453734
rect 380006 453498 380048 453734
rect 379728 453466 380048 453498
rect 410448 454054 410768 454086
rect 410448 453818 410490 454054
rect 410726 453818 410768 454054
rect 410448 453734 410768 453818
rect 410448 453498 410490 453734
rect 410726 453498 410768 453734
rect 410448 453466 410768 453498
rect 343888 450334 344208 450366
rect 343888 450098 343930 450334
rect 344166 450098 344208 450334
rect 343888 450014 344208 450098
rect 343888 449778 343930 450014
rect 344166 449778 344208 450014
rect 343888 449746 344208 449778
rect 374608 450334 374928 450366
rect 374608 450098 374650 450334
rect 374886 450098 374928 450334
rect 374608 450014 374928 450098
rect 374608 449778 374650 450014
rect 374886 449778 374928 450014
rect 374608 449746 374928 449778
rect 405328 450334 405648 450366
rect 405328 450098 405370 450334
rect 405606 450098 405648 450334
rect 405328 450014 405648 450098
rect 405328 449778 405370 450014
rect 405606 449778 405648 450014
rect 405328 449746 405648 449778
rect 338768 446614 339088 446646
rect 338768 446378 338810 446614
rect 339046 446378 339088 446614
rect 338768 446294 339088 446378
rect 338768 446058 338810 446294
rect 339046 446058 339088 446294
rect 338768 446026 339088 446058
rect 369488 446614 369808 446646
rect 369488 446378 369530 446614
rect 369766 446378 369808 446614
rect 369488 446294 369808 446378
rect 369488 446058 369530 446294
rect 369766 446058 369808 446294
rect 369488 446026 369808 446058
rect 400208 446614 400528 446646
rect 400208 446378 400250 446614
rect 400486 446378 400528 446614
rect 400208 446294 400528 446378
rect 400208 446058 400250 446294
rect 400486 446058 400528 446294
rect 400208 446026 400528 446058
rect 333648 442894 333968 442926
rect 333648 442658 333690 442894
rect 333926 442658 333968 442894
rect 333648 442574 333968 442658
rect 333648 442338 333690 442574
rect 333926 442338 333968 442574
rect 333648 442306 333968 442338
rect 364368 442894 364688 442926
rect 364368 442658 364410 442894
rect 364646 442658 364688 442894
rect 364368 442574 364688 442658
rect 364368 442338 364410 442574
rect 364646 442338 364688 442574
rect 364368 442306 364688 442338
rect 395088 442894 395408 442926
rect 395088 442658 395130 442894
rect 395366 442658 395408 442894
rect 395088 442574 395408 442658
rect 395088 442338 395130 442574
rect 395366 442338 395408 442574
rect 395088 442306 395408 442338
rect 328528 439174 328848 439206
rect 328528 438938 328570 439174
rect 328806 438938 328848 439174
rect 328528 438854 328848 438938
rect 328528 438618 328570 438854
rect 328806 438618 328848 438854
rect 328528 438586 328848 438618
rect 359248 439174 359568 439206
rect 359248 438938 359290 439174
rect 359526 438938 359568 439174
rect 359248 438854 359568 438938
rect 359248 438618 359290 438854
rect 359526 438618 359568 438854
rect 359248 438586 359568 438618
rect 389968 439174 390288 439206
rect 389968 438938 390010 439174
rect 390246 438938 390288 439174
rect 389968 438854 390288 438938
rect 389968 438618 390010 438854
rect 390246 438618 390288 438854
rect 389968 438586 390288 438618
rect 420688 439174 421008 439206
rect 420688 438938 420730 439174
rect 420966 438938 421008 439174
rect 420688 438854 421008 438938
rect 420688 438618 420730 438854
rect 420966 438618 421008 438854
rect 420688 438586 421008 438618
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 315834 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 316454 425494
rect 315834 425174 316454 425258
rect 315834 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 316454 425174
rect 313168 414334 313488 414366
rect 313168 414098 313210 414334
rect 313446 414098 313488 414334
rect 313168 414014 313488 414098
rect 313168 413778 313210 414014
rect 313446 413778 313488 414014
rect 313168 413746 313488 413778
rect 312114 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 312734 385774
rect 312114 385454 312734 385538
rect 312114 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 312734 385454
rect 308048 374614 308368 374646
rect 308048 374378 308090 374614
rect 308326 374378 308368 374614
rect 308048 374294 308368 374378
rect 308048 374058 308090 374294
rect 308326 374058 308368 374294
rect 308048 374026 308368 374058
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 302928 334894 303248 334926
rect 302928 334658 302970 334894
rect 303206 334658 303248 334894
rect 302928 334574 303248 334658
rect 302928 334338 302970 334574
rect 303206 334338 303248 334574
rect 302928 334306 303248 334338
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 287568 274054 287888 274086
rect 287568 273818 287610 274054
rect 287846 273818 287888 274054
rect 287568 273734 287888 273818
rect 287568 273498 287610 273734
rect 287846 273498 287888 273734
rect 287568 273466 287888 273498
rect 282448 270334 282768 270366
rect 282448 270098 282490 270334
rect 282726 270098 282768 270334
rect 282448 270014 282768 270098
rect 282448 269778 282490 270014
rect 282726 269778 282768 270014
rect 282448 269746 282768 269778
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 277328 230614 277648 230646
rect 277328 230378 277370 230614
rect 277606 230378 277648 230614
rect 277328 230294 277648 230378
rect 277328 230058 277370 230294
rect 277606 230058 277648 230294
rect 277328 230026 277648 230058
rect 276114 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 276734 205774
rect 276114 205454 276734 205538
rect 276114 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 276734 205454
rect 272208 190894 272528 190926
rect 272208 190658 272250 190894
rect 272486 190658 272528 190894
rect 272208 190574 272528 190658
rect 272208 190338 272250 190574
rect 272486 190338 272528 190574
rect 272208 190306 272528 190338
rect 268674 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 269294 162334
rect 268674 162014 269294 162098
rect 268674 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 269294 162014
rect 267088 151174 267408 151206
rect 267088 150938 267130 151174
rect 267366 150938 267408 151174
rect 267088 150854 267408 150938
rect 267088 150618 267130 150854
rect 267366 150618 267408 150854
rect 267088 150586 267408 150618
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 261968 111454 262288 111486
rect 261968 111218 262010 111454
rect 262246 111218 262288 111454
rect 261968 111134 262288 111218
rect 261968 110898 262010 111134
rect 262246 110898 262288 111134
rect 261968 110866 262288 110898
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 256848 58054 257168 58086
rect 256848 57818 256890 58054
rect 257126 57818 257168 58054
rect 256848 57734 257168 57818
rect 256848 57498 256890 57734
rect 257126 57498 257168 57734
rect 256848 57466 257168 57498
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 251728 18334 252048 18366
rect 251728 18098 251770 18334
rect 252006 18098 252048 18334
rect 251728 18014 252048 18098
rect 251728 17778 251770 18014
rect 252006 17778 252048 18014
rect 251728 17746 252048 17778
rect 246608 14614 246928 14646
rect 246608 14378 246650 14614
rect 246886 14378 246928 14614
rect 246608 14294 246928 14378
rect 246608 14058 246650 14294
rect 246886 14058 246928 14294
rect 246608 14026 246928 14058
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 3454 254414 38898
rect 257514 43174 258134 78618
rect 264954 86614 265574 122058
rect 268674 126334 269294 161778
rect 276114 169774 276734 205218
rect 279834 209494 280454 244938
rect 289794 255454 290414 290898
rect 292688 291454 293008 291486
rect 292688 291218 292730 291454
rect 292966 291218 293008 291454
rect 292688 291134 293008 291218
rect 292688 290898 292730 291134
rect 292966 290898 293008 291134
rect 292688 290866 293008 290898
rect 293514 259174 294134 294618
rect 297808 295174 298128 295206
rect 297808 294938 297850 295174
rect 298086 294938 298128 295174
rect 297808 294854 298128 294938
rect 297808 294618 297850 294854
rect 298086 294618 298128 294854
rect 297808 294586 298128 294618
rect 300954 266614 301574 302058
rect 304674 306334 305294 341778
rect 312114 349774 312734 385218
rect 315834 389494 316454 424938
rect 318288 418054 318608 418086
rect 318288 417818 318330 418054
rect 318566 417818 318608 418054
rect 318288 417734 318608 417818
rect 318288 417498 318330 417734
rect 318566 417498 318608 417734
rect 318288 417466 318608 417498
rect 323408 399454 323728 399486
rect 323408 399218 323450 399454
rect 323686 399218 323728 399454
rect 323408 399134 323728 399218
rect 323408 398898 323450 399134
rect 323686 398898 323728 399134
rect 323408 398866 323728 398898
rect 325794 399454 326414 434898
rect 354128 435454 354448 435486
rect 354128 435218 354170 435454
rect 354406 435218 354448 435454
rect 354128 435134 354448 435218
rect 354128 434898 354170 435134
rect 354406 434898 354448 435134
rect 354128 434866 354448 434898
rect 384848 435454 385168 435486
rect 384848 435218 384890 435454
rect 385126 435218 385168 435454
rect 384848 435134 385168 435218
rect 384848 434898 384890 435134
rect 385126 434898 385168 435134
rect 384848 434866 385168 434898
rect 415568 435454 415888 435486
rect 415568 435218 415610 435454
rect 415846 435218 415888 435454
rect 415568 435134 415888 435218
rect 415568 434898 415610 435134
rect 415846 434898 415888 435134
rect 415568 434866 415888 434898
rect 423834 425494 424454 460938
rect 433794 471454 434414 506898
rect 437514 511174 438134 546618
rect 444954 554614 445574 590058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 446288 579454 446608 579486
rect 446288 579218 446330 579454
rect 446566 579218 446608 579454
rect 446288 579134 446608 579218
rect 446288 578898 446330 579134
rect 446566 578898 446608 579134
rect 446288 578866 446608 578898
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 441168 526054 441488 526086
rect 441168 525818 441210 526054
rect 441446 525818 441488 526054
rect 441168 525734 441488 525818
rect 441168 525498 441210 525734
rect 441446 525498 441488 525734
rect 441168 525466 441488 525498
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 436048 486334 436368 486366
rect 436048 486098 436090 486334
rect 436326 486098 436368 486334
rect 436048 486014 436368 486098
rect 436048 485778 436090 486014
rect 436326 485778 436368 486014
rect 436048 485746 436368 485778
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 430928 446614 431248 446646
rect 430928 446378 430970 446614
rect 431206 446378 431248 446614
rect 430928 446294 431248 446378
rect 430928 446058 430970 446294
rect 431206 446058 431248 446294
rect 430928 446026 431248 446058
rect 425808 442894 426128 442926
rect 425808 442658 425850 442894
rect 426086 442658 426128 442894
rect 425808 442574 426128 442658
rect 425808 442338 425850 442574
rect 426086 442338 426128 442574
rect 425808 442306 426128 442338
rect 423834 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 424454 425494
rect 423834 425174 424454 425258
rect 423834 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 424454 425174
rect 349008 418054 349328 418086
rect 349008 417818 349050 418054
rect 349286 417818 349328 418054
rect 349008 417734 349328 417818
rect 349008 417498 349050 417734
rect 349286 417498 349328 417734
rect 349008 417466 349328 417498
rect 379728 418054 380048 418086
rect 379728 417818 379770 418054
rect 380006 417818 380048 418054
rect 379728 417734 380048 417818
rect 379728 417498 379770 417734
rect 380006 417498 380048 417734
rect 379728 417466 380048 417498
rect 410448 418054 410768 418086
rect 410448 417818 410490 418054
rect 410726 417818 410768 418054
rect 410448 417734 410768 417818
rect 410448 417498 410490 417734
rect 410726 417498 410768 417734
rect 410448 417466 410768 417498
rect 343888 414334 344208 414366
rect 343888 414098 343930 414334
rect 344166 414098 344208 414334
rect 343888 414014 344208 414098
rect 343888 413778 343930 414014
rect 344166 413778 344208 414014
rect 343888 413746 344208 413778
rect 374608 414334 374928 414366
rect 374608 414098 374650 414334
rect 374886 414098 374928 414334
rect 374608 414014 374928 414098
rect 374608 413778 374650 414014
rect 374886 413778 374928 414014
rect 374608 413746 374928 413778
rect 405328 414334 405648 414366
rect 405328 414098 405370 414334
rect 405606 414098 405648 414334
rect 405328 414014 405648 414098
rect 405328 413778 405370 414014
rect 405606 413778 405648 414014
rect 405328 413746 405648 413778
rect 338768 410614 339088 410646
rect 338768 410378 338810 410614
rect 339046 410378 339088 410614
rect 338768 410294 339088 410378
rect 338768 410058 338810 410294
rect 339046 410058 339088 410294
rect 338768 410026 339088 410058
rect 369488 410614 369808 410646
rect 369488 410378 369530 410614
rect 369766 410378 369808 410614
rect 369488 410294 369808 410378
rect 369488 410058 369530 410294
rect 369766 410058 369808 410294
rect 369488 410026 369808 410058
rect 400208 410614 400528 410646
rect 400208 410378 400250 410614
rect 400486 410378 400528 410614
rect 400208 410294 400528 410378
rect 400208 410058 400250 410294
rect 400486 410058 400528 410294
rect 400208 410026 400528 410058
rect 333648 406894 333968 406926
rect 333648 406658 333690 406894
rect 333926 406658 333968 406894
rect 333648 406574 333968 406658
rect 333648 406338 333690 406574
rect 333926 406338 333968 406574
rect 333648 406306 333968 406338
rect 364368 406894 364688 406926
rect 364368 406658 364410 406894
rect 364646 406658 364688 406894
rect 364368 406574 364688 406658
rect 364368 406338 364410 406574
rect 364646 406338 364688 406574
rect 364368 406306 364688 406338
rect 395088 406894 395408 406926
rect 395088 406658 395130 406894
rect 395366 406658 395408 406894
rect 395088 406574 395408 406658
rect 395088 406338 395130 406574
rect 395366 406338 395408 406574
rect 395088 406306 395408 406338
rect 328528 403174 328848 403206
rect 328528 402938 328570 403174
rect 328806 402938 328848 403174
rect 328528 402854 328848 402938
rect 328528 402618 328570 402854
rect 328806 402618 328848 402854
rect 328528 402586 328848 402618
rect 359248 403174 359568 403206
rect 359248 402938 359290 403174
rect 359526 402938 359568 403174
rect 359248 402854 359568 402938
rect 359248 402618 359290 402854
rect 359526 402618 359568 402854
rect 359248 402586 359568 402618
rect 389968 403174 390288 403206
rect 389968 402938 390010 403174
rect 390246 402938 390288 403174
rect 389968 402854 390288 402938
rect 389968 402618 390010 402854
rect 390246 402618 390288 402854
rect 389968 402586 390288 402618
rect 420688 403174 421008 403206
rect 420688 402938 420730 403174
rect 420966 402938 421008 403174
rect 420688 402854 421008 402938
rect 420688 402618 420730 402854
rect 420966 402618 421008 402854
rect 420688 402586 421008 402618
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 315834 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 316454 389494
rect 315834 389174 316454 389258
rect 315834 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 316454 389174
rect 313168 378334 313488 378366
rect 313168 378098 313210 378334
rect 313446 378098 313488 378334
rect 313168 378014 313488 378098
rect 313168 377778 313210 378014
rect 313446 377778 313488 378014
rect 313168 377746 313488 377778
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 308048 338614 308368 338646
rect 308048 338378 308090 338614
rect 308326 338378 308368 338614
rect 308048 338294 308368 338378
rect 308048 338058 308090 338294
rect 308326 338058 308368 338294
rect 308048 338026 308368 338058
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 302928 298894 303248 298926
rect 302928 298658 302970 298894
rect 303206 298658 303248 298894
rect 302928 298574 303248 298658
rect 302928 298338 302970 298574
rect 303206 298338 303248 298574
rect 302928 298306 303248 298338
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 287568 238054 287888 238086
rect 287568 237818 287610 238054
rect 287846 237818 287888 238054
rect 287568 237734 287888 237818
rect 287568 237498 287610 237734
rect 287846 237498 287888 237734
rect 287568 237466 287888 237498
rect 282448 234334 282768 234366
rect 282448 234098 282490 234334
rect 282726 234098 282768 234334
rect 282448 234014 282768 234098
rect 282448 233778 282490 234014
rect 282726 233778 282768 234014
rect 282448 233746 282768 233778
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 277328 194614 277648 194646
rect 277328 194378 277370 194614
rect 277606 194378 277648 194614
rect 277328 194294 277648 194378
rect 277328 194058 277370 194294
rect 277606 194058 277648 194294
rect 277328 194026 277648 194058
rect 276114 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 276734 169774
rect 276114 169454 276734 169538
rect 276114 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 276734 169454
rect 272208 154894 272528 154926
rect 272208 154658 272250 154894
rect 272486 154658 272528 154894
rect 272208 154574 272528 154658
rect 272208 154338 272250 154574
rect 272486 154338 272528 154574
rect 272208 154306 272528 154338
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 267088 115174 267408 115206
rect 267088 114938 267130 115174
rect 267366 114938 267408 115174
rect 267088 114854 267408 114938
rect 267088 114618 267130 114854
rect 267366 114618 267408 114854
rect 267088 114586 267408 114618
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 261968 75454 262288 75486
rect 261968 75218 262010 75454
rect 262246 75218 262288 75454
rect 261968 75134 262288 75218
rect 261968 74898 262010 75134
rect 262246 74898 262288 75134
rect 261968 74866 262288 74898
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 256848 22054 257168 22086
rect 256848 21818 256890 22054
rect 257126 21818 257168 22054
rect 256848 21734 257168 21818
rect 256848 21498 256890 21734
rect 257126 21498 257168 21734
rect 256848 21466 257168 21498
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 7174 258134 42618
rect 264954 50614 265574 86058
rect 268674 90334 269294 125778
rect 276114 133774 276734 169218
rect 279834 173494 280454 208938
rect 289794 219454 290414 254898
rect 292688 255454 293008 255486
rect 292688 255218 292730 255454
rect 292966 255218 293008 255454
rect 292688 255134 293008 255218
rect 292688 254898 292730 255134
rect 292966 254898 293008 255134
rect 292688 254866 293008 254898
rect 293514 223174 294134 258618
rect 297808 259174 298128 259206
rect 297808 258938 297850 259174
rect 298086 258938 298128 259174
rect 297808 258854 298128 258938
rect 297808 258618 297850 258854
rect 298086 258618 298128 258854
rect 297808 258586 298128 258618
rect 300954 230614 301574 266058
rect 304674 270334 305294 305778
rect 312114 313774 312734 349218
rect 315834 353494 316454 388938
rect 318288 382054 318608 382086
rect 318288 381818 318330 382054
rect 318566 381818 318608 382054
rect 318288 381734 318608 381818
rect 318288 381498 318330 381734
rect 318566 381498 318608 381734
rect 318288 381466 318608 381498
rect 323408 363454 323728 363486
rect 323408 363218 323450 363454
rect 323686 363218 323728 363454
rect 323408 363134 323728 363218
rect 323408 362898 323450 363134
rect 323686 362898 323728 363134
rect 323408 362866 323728 362898
rect 325794 363454 326414 398898
rect 354128 399454 354448 399486
rect 354128 399218 354170 399454
rect 354406 399218 354448 399454
rect 354128 399134 354448 399218
rect 354128 398898 354170 399134
rect 354406 398898 354448 399134
rect 354128 398866 354448 398898
rect 384848 399454 385168 399486
rect 384848 399218 384890 399454
rect 385126 399218 385168 399454
rect 384848 399134 385168 399218
rect 384848 398898 384890 399134
rect 385126 398898 385168 399134
rect 384848 398866 385168 398898
rect 415568 399454 415888 399486
rect 415568 399218 415610 399454
rect 415846 399218 415888 399454
rect 415568 399134 415888 399218
rect 415568 398898 415610 399134
rect 415846 398898 415888 399134
rect 415568 398866 415888 398898
rect 423834 389494 424454 424938
rect 433794 435454 434414 470898
rect 437514 475174 438134 510618
rect 444954 518614 445574 554058
rect 448674 558334 449294 593778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 602500 456734 637218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 451408 583174 451728 583206
rect 451408 582938 451450 583174
rect 451686 582938 451728 583174
rect 451408 582854 451728 582938
rect 451408 582618 451450 582854
rect 451686 582618 451728 582854
rect 451408 582586 451728 582618
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 446288 543454 446608 543486
rect 446288 543218 446330 543454
rect 446566 543218 446608 543454
rect 446288 543134 446608 543218
rect 446288 542898 446330 543134
rect 446566 542898 446608 543134
rect 446288 542866 446608 542898
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 441168 490054 441488 490086
rect 441168 489818 441210 490054
rect 441446 489818 441488 490054
rect 441168 489734 441488 489818
rect 441168 489498 441210 489734
rect 441446 489498 441488 489734
rect 441168 489466 441488 489498
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 436048 450334 436368 450366
rect 436048 450098 436090 450334
rect 436326 450098 436368 450334
rect 436048 450014 436368 450098
rect 436048 449778 436090 450014
rect 436326 449778 436368 450014
rect 436048 449746 436368 449778
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 430928 410614 431248 410646
rect 430928 410378 430970 410614
rect 431206 410378 431248 410614
rect 430928 410294 431248 410378
rect 430928 410058 430970 410294
rect 431206 410058 431248 410294
rect 430928 410026 431248 410058
rect 425808 406894 426128 406926
rect 425808 406658 425850 406894
rect 426086 406658 426128 406894
rect 425808 406574 426128 406658
rect 425808 406338 425850 406574
rect 426086 406338 426128 406574
rect 425808 406306 426128 406338
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 349008 382054 349328 382086
rect 349008 381818 349050 382054
rect 349286 381818 349328 382054
rect 349008 381734 349328 381818
rect 349008 381498 349050 381734
rect 349286 381498 349328 381734
rect 349008 381466 349328 381498
rect 379728 382054 380048 382086
rect 379728 381818 379770 382054
rect 380006 381818 380048 382054
rect 379728 381734 380048 381818
rect 379728 381498 379770 381734
rect 380006 381498 380048 381734
rect 379728 381466 380048 381498
rect 410448 382054 410768 382086
rect 410448 381818 410490 382054
rect 410726 381818 410768 382054
rect 410448 381734 410768 381818
rect 410448 381498 410490 381734
rect 410726 381498 410768 381734
rect 410448 381466 410768 381498
rect 343888 378334 344208 378366
rect 343888 378098 343930 378334
rect 344166 378098 344208 378334
rect 343888 378014 344208 378098
rect 343888 377778 343930 378014
rect 344166 377778 344208 378014
rect 343888 377746 344208 377778
rect 374608 378334 374928 378366
rect 374608 378098 374650 378334
rect 374886 378098 374928 378334
rect 374608 378014 374928 378098
rect 374608 377778 374650 378014
rect 374886 377778 374928 378014
rect 374608 377746 374928 377778
rect 405328 378334 405648 378366
rect 405328 378098 405370 378334
rect 405606 378098 405648 378334
rect 405328 378014 405648 378098
rect 405328 377778 405370 378014
rect 405606 377778 405648 378014
rect 405328 377746 405648 377778
rect 338768 374614 339088 374646
rect 338768 374378 338810 374614
rect 339046 374378 339088 374614
rect 338768 374294 339088 374378
rect 338768 374058 338810 374294
rect 339046 374058 339088 374294
rect 338768 374026 339088 374058
rect 369488 374614 369808 374646
rect 369488 374378 369530 374614
rect 369766 374378 369808 374614
rect 369488 374294 369808 374378
rect 369488 374058 369530 374294
rect 369766 374058 369808 374294
rect 369488 374026 369808 374058
rect 400208 374614 400528 374646
rect 400208 374378 400250 374614
rect 400486 374378 400528 374614
rect 400208 374294 400528 374378
rect 400208 374058 400250 374294
rect 400486 374058 400528 374294
rect 400208 374026 400528 374058
rect 333648 370894 333968 370926
rect 333648 370658 333690 370894
rect 333926 370658 333968 370894
rect 333648 370574 333968 370658
rect 333648 370338 333690 370574
rect 333926 370338 333968 370574
rect 333648 370306 333968 370338
rect 364368 370894 364688 370926
rect 364368 370658 364410 370894
rect 364646 370658 364688 370894
rect 364368 370574 364688 370658
rect 364368 370338 364410 370574
rect 364646 370338 364688 370574
rect 364368 370306 364688 370338
rect 395088 370894 395408 370926
rect 395088 370658 395130 370894
rect 395366 370658 395408 370894
rect 395088 370574 395408 370658
rect 395088 370338 395130 370574
rect 395366 370338 395408 370574
rect 395088 370306 395408 370338
rect 328528 367174 328848 367206
rect 328528 366938 328570 367174
rect 328806 366938 328848 367174
rect 328528 366854 328848 366938
rect 328528 366618 328570 366854
rect 328806 366618 328848 366854
rect 328528 366586 328848 366618
rect 359248 367174 359568 367206
rect 359248 366938 359290 367174
rect 359526 366938 359568 367174
rect 359248 366854 359568 366938
rect 359248 366618 359290 366854
rect 359526 366618 359568 366854
rect 359248 366586 359568 366618
rect 389968 367174 390288 367206
rect 389968 366938 390010 367174
rect 390246 366938 390288 367174
rect 389968 366854 390288 366938
rect 389968 366618 390010 366854
rect 390246 366618 390288 366854
rect 389968 366586 390288 366618
rect 420688 367174 421008 367206
rect 420688 366938 420730 367174
rect 420966 366938 421008 367174
rect 420688 366854 421008 366938
rect 420688 366618 420730 366854
rect 420966 366618 421008 366854
rect 420688 366586 421008 366618
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 313168 342334 313488 342366
rect 313168 342098 313210 342334
rect 313446 342098 313488 342334
rect 313168 342014 313488 342098
rect 313168 341778 313210 342014
rect 313446 341778 313488 342014
rect 313168 341746 313488 341778
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 308048 302614 308368 302646
rect 308048 302378 308090 302614
rect 308326 302378 308368 302614
rect 308048 302294 308368 302378
rect 308048 302058 308090 302294
rect 308326 302058 308368 302294
rect 308048 302026 308368 302058
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 302928 262894 303248 262926
rect 302928 262658 302970 262894
rect 303206 262658 303248 262894
rect 302928 262574 303248 262658
rect 302928 262338 302970 262574
rect 303206 262338 303248 262574
rect 302928 262306 303248 262338
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 287568 202054 287888 202086
rect 287568 201818 287610 202054
rect 287846 201818 287888 202054
rect 287568 201734 287888 201818
rect 287568 201498 287610 201734
rect 287846 201498 287888 201734
rect 287568 201466 287888 201498
rect 282448 198334 282768 198366
rect 282448 198098 282490 198334
rect 282726 198098 282768 198334
rect 282448 198014 282768 198098
rect 282448 197778 282490 198014
rect 282726 197778 282768 198014
rect 282448 197746 282768 197778
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 277328 158614 277648 158646
rect 277328 158378 277370 158614
rect 277606 158378 277648 158614
rect 277328 158294 277648 158378
rect 277328 158058 277370 158294
rect 277606 158058 277648 158294
rect 277328 158026 277648 158058
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 272208 118894 272528 118926
rect 272208 118658 272250 118894
rect 272486 118658 272528 118894
rect 272208 118574 272528 118658
rect 272208 118338 272250 118574
rect 272486 118338 272528 118574
rect 272208 118306 272528 118338
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 267088 79174 267408 79206
rect 267088 78938 267130 79174
rect 267366 78938 267408 79174
rect 267088 78854 267408 78938
rect 267088 78618 267130 78854
rect 267366 78618 267408 78854
rect 267088 78586 267408 78618
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 261968 39454 262288 39486
rect 261968 39218 262010 39454
rect 262246 39218 262288 39454
rect 261968 39134 262288 39218
rect 261968 38898 262010 39134
rect 262246 38898 262288 39134
rect 261968 38866 262288 38898
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 264954 14614 265574 50058
rect 268674 54334 269294 89778
rect 276114 97774 276734 133218
rect 279834 137494 280454 172938
rect 289794 183454 290414 218898
rect 292688 219454 293008 219486
rect 292688 219218 292730 219454
rect 292966 219218 293008 219454
rect 292688 219134 293008 219218
rect 292688 218898 292730 219134
rect 292966 218898 293008 219134
rect 292688 218866 293008 218898
rect 293514 187174 294134 222618
rect 297808 223174 298128 223206
rect 297808 222938 297850 223174
rect 298086 222938 298128 223174
rect 297808 222854 298128 222938
rect 297808 222618 297850 222854
rect 298086 222618 298128 222854
rect 297808 222586 298128 222618
rect 300954 194614 301574 230058
rect 304674 234334 305294 269778
rect 312114 277774 312734 313218
rect 315834 317494 316454 352938
rect 318288 346054 318608 346086
rect 318288 345818 318330 346054
rect 318566 345818 318608 346054
rect 318288 345734 318608 345818
rect 318288 345498 318330 345734
rect 318566 345498 318608 345734
rect 318288 345466 318608 345498
rect 323408 327454 323728 327486
rect 323408 327218 323450 327454
rect 323686 327218 323728 327454
rect 323408 327134 323728 327218
rect 323408 326898 323450 327134
rect 323686 326898 323728 327134
rect 323408 326866 323728 326898
rect 325794 327454 326414 362898
rect 354128 363454 354448 363486
rect 354128 363218 354170 363454
rect 354406 363218 354448 363454
rect 354128 363134 354448 363218
rect 354128 362898 354170 363134
rect 354406 362898 354448 363134
rect 354128 362866 354448 362898
rect 384848 363454 385168 363486
rect 384848 363218 384890 363454
rect 385126 363218 385168 363454
rect 384848 363134 385168 363218
rect 384848 362898 384890 363134
rect 385126 362898 385168 363134
rect 384848 362866 385168 362898
rect 415568 363454 415888 363486
rect 415568 363218 415610 363454
rect 415846 363218 415888 363454
rect 415568 363134 415888 363218
rect 415568 362898 415610 363134
rect 415846 362898 415888 363134
rect 415568 362866 415888 362898
rect 423834 353494 424454 388938
rect 433794 399454 434414 434898
rect 437514 439174 438134 474618
rect 444954 482614 445574 518058
rect 448674 522334 449294 557778
rect 452394 562054 453014 597498
rect 456528 586894 456848 586926
rect 456528 586658 456570 586894
rect 456806 586658 456848 586894
rect 456528 586574 456848 586658
rect 456528 586338 456570 586574
rect 456806 586338 456848 586574
rect 456528 586306 456848 586338
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 451408 547174 451728 547206
rect 451408 546938 451450 547174
rect 451686 546938 451728 547174
rect 451408 546854 451728 546938
rect 451408 546618 451450 546854
rect 451686 546618 451728 546854
rect 451408 546586 451728 546618
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 446288 507454 446608 507486
rect 446288 507218 446330 507454
rect 446566 507218 446608 507454
rect 446288 507134 446608 507218
rect 446288 506898 446330 507134
rect 446566 506898 446608 507134
rect 446288 506866 446608 506898
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 441168 454054 441488 454086
rect 441168 453818 441210 454054
rect 441446 453818 441488 454054
rect 441168 453734 441488 453818
rect 441168 453498 441210 453734
rect 441446 453498 441488 453734
rect 441168 453466 441488 453498
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 436048 414334 436368 414366
rect 436048 414098 436090 414334
rect 436326 414098 436368 414334
rect 436048 414014 436368 414098
rect 436048 413778 436090 414014
rect 436326 413778 436368 414014
rect 436048 413746 436368 413778
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 430928 374614 431248 374646
rect 430928 374378 430970 374614
rect 431206 374378 431248 374614
rect 430928 374294 431248 374378
rect 430928 374058 430970 374294
rect 431206 374058 431248 374294
rect 430928 374026 431248 374058
rect 425808 370894 426128 370926
rect 425808 370658 425850 370894
rect 426086 370658 426128 370894
rect 425808 370574 426128 370658
rect 425808 370338 425850 370574
rect 426086 370338 426128 370574
rect 425808 370306 426128 370338
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 349008 346054 349328 346086
rect 349008 345818 349050 346054
rect 349286 345818 349328 346054
rect 349008 345734 349328 345818
rect 349008 345498 349050 345734
rect 349286 345498 349328 345734
rect 349008 345466 349328 345498
rect 379728 346054 380048 346086
rect 379728 345818 379770 346054
rect 380006 345818 380048 346054
rect 379728 345734 380048 345818
rect 379728 345498 379770 345734
rect 380006 345498 380048 345734
rect 379728 345466 380048 345498
rect 410448 346054 410768 346086
rect 410448 345818 410490 346054
rect 410726 345818 410768 346054
rect 410448 345734 410768 345818
rect 410448 345498 410490 345734
rect 410726 345498 410768 345734
rect 410448 345466 410768 345498
rect 343888 342334 344208 342366
rect 343888 342098 343930 342334
rect 344166 342098 344208 342334
rect 343888 342014 344208 342098
rect 343888 341778 343930 342014
rect 344166 341778 344208 342014
rect 343888 341746 344208 341778
rect 374608 342334 374928 342366
rect 374608 342098 374650 342334
rect 374886 342098 374928 342334
rect 374608 342014 374928 342098
rect 374608 341778 374650 342014
rect 374886 341778 374928 342014
rect 374608 341746 374928 341778
rect 405328 342334 405648 342366
rect 405328 342098 405370 342334
rect 405606 342098 405648 342334
rect 405328 342014 405648 342098
rect 405328 341778 405370 342014
rect 405606 341778 405648 342014
rect 405328 341746 405648 341778
rect 338768 338614 339088 338646
rect 338768 338378 338810 338614
rect 339046 338378 339088 338614
rect 338768 338294 339088 338378
rect 338768 338058 338810 338294
rect 339046 338058 339088 338294
rect 338768 338026 339088 338058
rect 369488 338614 369808 338646
rect 369488 338378 369530 338614
rect 369766 338378 369808 338614
rect 369488 338294 369808 338378
rect 369488 338058 369530 338294
rect 369766 338058 369808 338294
rect 369488 338026 369808 338058
rect 400208 338614 400528 338646
rect 400208 338378 400250 338614
rect 400486 338378 400528 338614
rect 400208 338294 400528 338378
rect 400208 338058 400250 338294
rect 400486 338058 400528 338294
rect 400208 338026 400528 338058
rect 333648 334894 333968 334926
rect 333648 334658 333690 334894
rect 333926 334658 333968 334894
rect 333648 334574 333968 334658
rect 333648 334338 333690 334574
rect 333926 334338 333968 334574
rect 333648 334306 333968 334338
rect 364368 334894 364688 334926
rect 364368 334658 364410 334894
rect 364646 334658 364688 334894
rect 364368 334574 364688 334658
rect 364368 334338 364410 334574
rect 364646 334338 364688 334574
rect 364368 334306 364688 334338
rect 395088 334894 395408 334926
rect 395088 334658 395130 334894
rect 395366 334658 395408 334894
rect 395088 334574 395408 334658
rect 395088 334338 395130 334574
rect 395366 334338 395408 334574
rect 395088 334306 395408 334338
rect 328528 331174 328848 331206
rect 328528 330938 328570 331174
rect 328806 330938 328848 331174
rect 328528 330854 328848 330938
rect 328528 330618 328570 330854
rect 328806 330618 328848 330854
rect 328528 330586 328848 330618
rect 359248 331174 359568 331206
rect 359248 330938 359290 331174
rect 359526 330938 359568 331174
rect 359248 330854 359568 330938
rect 359248 330618 359290 330854
rect 359526 330618 359568 330854
rect 359248 330586 359568 330618
rect 389968 331174 390288 331206
rect 389968 330938 390010 331174
rect 390246 330938 390288 331174
rect 389968 330854 390288 330938
rect 389968 330618 390010 330854
rect 390246 330618 390288 330854
rect 389968 330586 390288 330618
rect 420688 331174 421008 331206
rect 420688 330938 420730 331174
rect 420966 330938 421008 331174
rect 420688 330854 421008 330938
rect 420688 330618 420730 330854
rect 420966 330618 421008 330854
rect 420688 330586 421008 330618
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 313168 306334 313488 306366
rect 313168 306098 313210 306334
rect 313446 306098 313488 306334
rect 313168 306014 313488 306098
rect 313168 305778 313210 306014
rect 313446 305778 313488 306014
rect 313168 305746 313488 305778
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 308048 266614 308368 266646
rect 308048 266378 308090 266614
rect 308326 266378 308368 266614
rect 308048 266294 308368 266378
rect 308048 266058 308090 266294
rect 308326 266058 308368 266294
rect 308048 266026 308368 266058
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 302928 226894 303248 226926
rect 302928 226658 302970 226894
rect 303206 226658 303248 226894
rect 302928 226574 303248 226658
rect 302928 226338 302970 226574
rect 303206 226338 303248 226574
rect 302928 226306 303248 226338
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 287568 166054 287888 166086
rect 287568 165818 287610 166054
rect 287846 165818 287888 166054
rect 287568 165734 287888 165818
rect 287568 165498 287610 165734
rect 287846 165498 287888 165734
rect 287568 165466 287888 165498
rect 282448 162334 282768 162366
rect 282448 162098 282490 162334
rect 282726 162098 282768 162334
rect 282448 162014 282768 162098
rect 282448 161778 282490 162014
rect 282726 161778 282768 162014
rect 282448 161746 282768 161778
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 277328 122614 277648 122646
rect 277328 122378 277370 122614
rect 277606 122378 277648 122614
rect 277328 122294 277648 122378
rect 277328 122058 277370 122294
rect 277606 122058 277648 122294
rect 277328 122026 277648 122058
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 272208 82894 272528 82926
rect 272208 82658 272250 82894
rect 272486 82658 272528 82894
rect 272208 82574 272528 82658
rect 272208 82338 272250 82574
rect 272486 82338 272528 82574
rect 272208 82306 272528 82338
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 267088 43174 267408 43206
rect 267088 42938 267130 43174
rect 267366 42938 267408 43174
rect 267088 42854 267408 42938
rect 267088 42618 267130 42854
rect 267366 42618 267408 42854
rect 267088 42586 267408 42618
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 -2266 261854 2988
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 -3226 265574 14058
rect 268674 18334 269294 53778
rect 276114 61774 276734 97218
rect 279834 101494 280454 136938
rect 289794 147454 290414 182898
rect 292688 183454 293008 183486
rect 292688 183218 292730 183454
rect 292966 183218 293008 183454
rect 292688 183134 293008 183218
rect 292688 182898 292730 183134
rect 292966 182898 293008 183134
rect 292688 182866 293008 182898
rect 293514 151174 294134 186618
rect 297808 187174 298128 187206
rect 297808 186938 297850 187174
rect 298086 186938 298128 187174
rect 297808 186854 298128 186938
rect 297808 186618 297850 186854
rect 298086 186618 298128 186854
rect 297808 186586 298128 186618
rect 300954 158614 301574 194058
rect 304674 198334 305294 233778
rect 312114 241774 312734 277218
rect 315834 281494 316454 316938
rect 318288 310054 318608 310086
rect 318288 309818 318330 310054
rect 318566 309818 318608 310054
rect 318288 309734 318608 309818
rect 318288 309498 318330 309734
rect 318566 309498 318608 309734
rect 318288 309466 318608 309498
rect 323408 291454 323728 291486
rect 323408 291218 323450 291454
rect 323686 291218 323728 291454
rect 323408 291134 323728 291218
rect 323408 290898 323450 291134
rect 323686 290898 323728 291134
rect 323408 290866 323728 290898
rect 325794 291454 326414 326898
rect 354128 327454 354448 327486
rect 354128 327218 354170 327454
rect 354406 327218 354448 327454
rect 354128 327134 354448 327218
rect 354128 326898 354170 327134
rect 354406 326898 354448 327134
rect 354128 326866 354448 326898
rect 384848 327454 385168 327486
rect 384848 327218 384890 327454
rect 385126 327218 385168 327454
rect 384848 327134 385168 327218
rect 384848 326898 384890 327134
rect 385126 326898 385168 327134
rect 384848 326866 385168 326898
rect 415568 327454 415888 327486
rect 415568 327218 415610 327454
rect 415846 327218 415888 327454
rect 415568 327134 415888 327218
rect 415568 326898 415610 327134
rect 415846 326898 415888 327134
rect 415568 326866 415888 326898
rect 423834 317494 424454 352938
rect 433794 363454 434414 398898
rect 437514 403174 438134 438618
rect 444954 446614 445574 482058
rect 448674 486334 449294 521778
rect 452394 526054 453014 561498
rect 459834 569494 460454 604938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 466768 594334 467088 594366
rect 466768 594098 466810 594334
rect 467046 594098 467088 594334
rect 466768 594014 467088 594098
rect 466768 593778 466810 594014
rect 467046 593778 467088 594014
rect 466768 593746 467088 593778
rect 461648 590614 461968 590646
rect 461648 590378 461690 590614
rect 461926 590378 461968 590614
rect 461648 590294 461968 590378
rect 461648 590058 461690 590294
rect 461926 590058 461968 590294
rect 461648 590026 461968 590058
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 456528 550894 456848 550926
rect 456528 550658 456570 550894
rect 456806 550658 456848 550894
rect 456528 550574 456848 550658
rect 456528 550338 456570 550574
rect 456806 550338 456848 550574
rect 456528 550306 456848 550338
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 451408 511174 451728 511206
rect 451408 510938 451450 511174
rect 451686 510938 451728 511174
rect 451408 510854 451728 510938
rect 451408 510618 451450 510854
rect 451686 510618 451728 510854
rect 451408 510586 451728 510618
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 446288 471454 446608 471486
rect 446288 471218 446330 471454
rect 446566 471218 446608 471454
rect 446288 471134 446608 471218
rect 446288 470898 446330 471134
rect 446566 470898 446608 471134
rect 446288 470866 446608 470898
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 441168 418054 441488 418086
rect 441168 417818 441210 418054
rect 441446 417818 441488 418054
rect 441168 417734 441488 417818
rect 441168 417498 441210 417734
rect 441446 417498 441488 417734
rect 441168 417466 441488 417498
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 436048 378334 436368 378366
rect 436048 378098 436090 378334
rect 436326 378098 436368 378334
rect 436048 378014 436368 378098
rect 436048 377778 436090 378014
rect 436326 377778 436368 378014
rect 436048 377746 436368 377778
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 430928 338614 431248 338646
rect 430928 338378 430970 338614
rect 431206 338378 431248 338614
rect 430928 338294 431248 338378
rect 430928 338058 430970 338294
rect 431206 338058 431248 338294
rect 430928 338026 431248 338058
rect 425808 334894 426128 334926
rect 425808 334658 425850 334894
rect 426086 334658 426128 334894
rect 425808 334574 426128 334658
rect 425808 334338 425850 334574
rect 426086 334338 426128 334574
rect 425808 334306 426128 334338
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 349008 310054 349328 310086
rect 349008 309818 349050 310054
rect 349286 309818 349328 310054
rect 349008 309734 349328 309818
rect 349008 309498 349050 309734
rect 349286 309498 349328 309734
rect 349008 309466 349328 309498
rect 379728 310054 380048 310086
rect 379728 309818 379770 310054
rect 380006 309818 380048 310054
rect 379728 309734 380048 309818
rect 379728 309498 379770 309734
rect 380006 309498 380048 309734
rect 379728 309466 380048 309498
rect 410448 310054 410768 310086
rect 410448 309818 410490 310054
rect 410726 309818 410768 310054
rect 410448 309734 410768 309818
rect 410448 309498 410490 309734
rect 410726 309498 410768 309734
rect 410448 309466 410768 309498
rect 343888 306334 344208 306366
rect 343888 306098 343930 306334
rect 344166 306098 344208 306334
rect 343888 306014 344208 306098
rect 343888 305778 343930 306014
rect 344166 305778 344208 306014
rect 343888 305746 344208 305778
rect 374608 306334 374928 306366
rect 374608 306098 374650 306334
rect 374886 306098 374928 306334
rect 374608 306014 374928 306098
rect 374608 305778 374650 306014
rect 374886 305778 374928 306014
rect 374608 305746 374928 305778
rect 405328 306334 405648 306366
rect 405328 306098 405370 306334
rect 405606 306098 405648 306334
rect 405328 306014 405648 306098
rect 405328 305778 405370 306014
rect 405606 305778 405648 306014
rect 405328 305746 405648 305778
rect 338768 302614 339088 302646
rect 338768 302378 338810 302614
rect 339046 302378 339088 302614
rect 338768 302294 339088 302378
rect 338768 302058 338810 302294
rect 339046 302058 339088 302294
rect 338768 302026 339088 302058
rect 369488 302614 369808 302646
rect 369488 302378 369530 302614
rect 369766 302378 369808 302614
rect 369488 302294 369808 302378
rect 369488 302058 369530 302294
rect 369766 302058 369808 302294
rect 369488 302026 369808 302058
rect 400208 302614 400528 302646
rect 400208 302378 400250 302614
rect 400486 302378 400528 302614
rect 400208 302294 400528 302378
rect 400208 302058 400250 302294
rect 400486 302058 400528 302294
rect 400208 302026 400528 302058
rect 333648 298894 333968 298926
rect 333648 298658 333690 298894
rect 333926 298658 333968 298894
rect 333648 298574 333968 298658
rect 333648 298338 333690 298574
rect 333926 298338 333968 298574
rect 333648 298306 333968 298338
rect 364368 298894 364688 298926
rect 364368 298658 364410 298894
rect 364646 298658 364688 298894
rect 364368 298574 364688 298658
rect 364368 298338 364410 298574
rect 364646 298338 364688 298574
rect 364368 298306 364688 298338
rect 395088 298894 395408 298926
rect 395088 298658 395130 298894
rect 395366 298658 395408 298894
rect 395088 298574 395408 298658
rect 395088 298338 395130 298574
rect 395366 298338 395408 298574
rect 395088 298306 395408 298338
rect 328528 295174 328848 295206
rect 328528 294938 328570 295174
rect 328806 294938 328848 295174
rect 328528 294854 328848 294938
rect 328528 294618 328570 294854
rect 328806 294618 328848 294854
rect 328528 294586 328848 294618
rect 359248 295174 359568 295206
rect 359248 294938 359290 295174
rect 359526 294938 359568 295174
rect 359248 294854 359568 294938
rect 359248 294618 359290 294854
rect 359526 294618 359568 294854
rect 359248 294586 359568 294618
rect 389968 295174 390288 295206
rect 389968 294938 390010 295174
rect 390246 294938 390288 295174
rect 389968 294854 390288 294938
rect 389968 294618 390010 294854
rect 390246 294618 390288 294854
rect 389968 294586 390288 294618
rect 420688 295174 421008 295206
rect 420688 294938 420730 295174
rect 420966 294938 421008 295174
rect 420688 294854 421008 294938
rect 420688 294618 420730 294854
rect 420966 294618 421008 294854
rect 420688 294586 421008 294618
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 313168 270334 313488 270366
rect 313168 270098 313210 270334
rect 313446 270098 313488 270334
rect 313168 270014 313488 270098
rect 313168 269778 313210 270014
rect 313446 269778 313488 270014
rect 313168 269746 313488 269778
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 308048 230614 308368 230646
rect 308048 230378 308090 230614
rect 308326 230378 308368 230614
rect 308048 230294 308368 230378
rect 308048 230058 308090 230294
rect 308326 230058 308368 230294
rect 308048 230026 308368 230058
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 302928 190894 303248 190926
rect 302928 190658 302970 190894
rect 303206 190658 303248 190894
rect 302928 190574 303248 190658
rect 302928 190338 302970 190574
rect 303206 190338 303248 190574
rect 302928 190306 303248 190338
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 287568 130054 287888 130086
rect 287568 129818 287610 130054
rect 287846 129818 287888 130054
rect 287568 129734 287888 129818
rect 287568 129498 287610 129734
rect 287846 129498 287888 129734
rect 287568 129466 287888 129498
rect 282448 126334 282768 126366
rect 282448 126098 282490 126334
rect 282726 126098 282768 126334
rect 282448 126014 282768 126098
rect 282448 125778 282490 126014
rect 282726 125778 282768 126014
rect 282448 125746 282768 125778
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 277328 86614 277648 86646
rect 277328 86378 277370 86614
rect 277606 86378 277648 86614
rect 277328 86294 277648 86378
rect 277328 86058 277370 86294
rect 277606 86058 277648 86294
rect 277328 86026 277648 86058
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 272208 46894 272528 46926
rect 272208 46658 272250 46894
rect 272486 46658 272528 46894
rect 272208 46574 272528 46658
rect 272208 46338 272250 46574
rect 272486 46338 272528 46574
rect 272208 46306 272528 46338
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 267088 7174 267408 7206
rect 267088 6938 267130 7174
rect 267366 6938 267408 7174
rect 267088 6854 267408 6938
rect 267088 6618 267130 6854
rect 267366 6618 267408 6854
rect 267088 6586 267408 6618
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 -4186 269294 17778
rect 276114 25774 276734 61218
rect 279834 65494 280454 100938
rect 289794 111454 290414 146898
rect 292688 147454 293008 147486
rect 292688 147218 292730 147454
rect 292966 147218 293008 147454
rect 292688 147134 293008 147218
rect 292688 146898 292730 147134
rect 292966 146898 293008 147134
rect 292688 146866 293008 146898
rect 293514 115174 294134 150618
rect 297808 151174 298128 151206
rect 297808 150938 297850 151174
rect 298086 150938 298128 151174
rect 297808 150854 298128 150938
rect 297808 150618 297850 150854
rect 298086 150618 298128 150854
rect 297808 150586 298128 150618
rect 300954 122614 301574 158058
rect 304674 162334 305294 197778
rect 312114 205774 312734 241218
rect 315834 245494 316454 280938
rect 318288 274054 318608 274086
rect 318288 273818 318330 274054
rect 318566 273818 318608 274054
rect 318288 273734 318608 273818
rect 318288 273498 318330 273734
rect 318566 273498 318608 273734
rect 318288 273466 318608 273498
rect 323408 255454 323728 255486
rect 323408 255218 323450 255454
rect 323686 255218 323728 255454
rect 323408 255134 323728 255218
rect 323408 254898 323450 255134
rect 323686 254898 323728 255134
rect 323408 254866 323728 254898
rect 325794 255454 326414 290898
rect 354128 291454 354448 291486
rect 354128 291218 354170 291454
rect 354406 291218 354448 291454
rect 354128 291134 354448 291218
rect 354128 290898 354170 291134
rect 354406 290898 354448 291134
rect 354128 290866 354448 290898
rect 384848 291454 385168 291486
rect 384848 291218 384890 291454
rect 385126 291218 385168 291454
rect 384848 291134 385168 291218
rect 384848 290898 384890 291134
rect 385126 290898 385168 291134
rect 384848 290866 385168 290898
rect 415568 291454 415888 291486
rect 415568 291218 415610 291454
rect 415846 291218 415888 291454
rect 415568 291134 415888 291218
rect 415568 290898 415610 291134
rect 415846 290898 415888 291134
rect 415568 290866 415888 290898
rect 423834 281494 424454 316938
rect 433794 327454 434414 362898
rect 437514 367174 438134 402618
rect 444954 410614 445574 446058
rect 448674 450334 449294 485778
rect 452394 490054 453014 525498
rect 459834 533494 460454 568938
rect 469794 579454 470414 614898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 471888 598054 472208 598086
rect 471888 597818 471930 598054
rect 472166 597818 472208 598054
rect 471888 597734 472208 597818
rect 471888 597498 471930 597734
rect 472166 597498 472208 597734
rect 471888 597466 472208 597498
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 466768 558334 467088 558366
rect 466768 558098 466810 558334
rect 467046 558098 467088 558334
rect 466768 558014 467088 558098
rect 466768 557778 466810 558014
rect 467046 557778 467088 558014
rect 466768 557746 467088 557778
rect 461648 554614 461968 554646
rect 461648 554378 461690 554614
rect 461926 554378 461968 554614
rect 461648 554294 461968 554378
rect 461648 554058 461690 554294
rect 461926 554058 461968 554294
rect 461648 554026 461968 554058
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 456528 514894 456848 514926
rect 456528 514658 456570 514894
rect 456806 514658 456848 514894
rect 456528 514574 456848 514658
rect 456528 514338 456570 514574
rect 456806 514338 456848 514574
rect 456528 514306 456848 514338
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 451408 475174 451728 475206
rect 451408 474938 451450 475174
rect 451686 474938 451728 475174
rect 451408 474854 451728 474938
rect 451408 474618 451450 474854
rect 451686 474618 451728 474854
rect 451408 474586 451728 474618
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 446288 435454 446608 435486
rect 446288 435218 446330 435454
rect 446566 435218 446608 435454
rect 446288 435134 446608 435218
rect 446288 434898 446330 435134
rect 446566 434898 446608 435134
rect 446288 434866 446608 434898
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 441168 382054 441488 382086
rect 441168 381818 441210 382054
rect 441446 381818 441488 382054
rect 441168 381734 441488 381818
rect 441168 381498 441210 381734
rect 441446 381498 441488 381734
rect 441168 381466 441488 381498
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 436048 342334 436368 342366
rect 436048 342098 436090 342334
rect 436326 342098 436368 342334
rect 436048 342014 436368 342098
rect 436048 341778 436090 342014
rect 436326 341778 436368 342014
rect 436048 341746 436368 341778
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 430928 302614 431248 302646
rect 430928 302378 430970 302614
rect 431206 302378 431248 302614
rect 430928 302294 431248 302378
rect 430928 302058 430970 302294
rect 431206 302058 431248 302294
rect 430928 302026 431248 302058
rect 425808 298894 426128 298926
rect 425808 298658 425850 298894
rect 426086 298658 426128 298894
rect 425808 298574 426128 298658
rect 425808 298338 425850 298574
rect 426086 298338 426128 298574
rect 425808 298306 426128 298338
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 349008 274054 349328 274086
rect 349008 273818 349050 274054
rect 349286 273818 349328 274054
rect 349008 273734 349328 273818
rect 349008 273498 349050 273734
rect 349286 273498 349328 273734
rect 349008 273466 349328 273498
rect 379728 274054 380048 274086
rect 379728 273818 379770 274054
rect 380006 273818 380048 274054
rect 379728 273734 380048 273818
rect 379728 273498 379770 273734
rect 380006 273498 380048 273734
rect 379728 273466 380048 273498
rect 410448 274054 410768 274086
rect 410448 273818 410490 274054
rect 410726 273818 410768 274054
rect 410448 273734 410768 273818
rect 410448 273498 410490 273734
rect 410726 273498 410768 273734
rect 410448 273466 410768 273498
rect 343888 270334 344208 270366
rect 343888 270098 343930 270334
rect 344166 270098 344208 270334
rect 343888 270014 344208 270098
rect 343888 269778 343930 270014
rect 344166 269778 344208 270014
rect 343888 269746 344208 269778
rect 374608 270334 374928 270366
rect 374608 270098 374650 270334
rect 374886 270098 374928 270334
rect 374608 270014 374928 270098
rect 374608 269778 374650 270014
rect 374886 269778 374928 270014
rect 374608 269746 374928 269778
rect 405328 270334 405648 270366
rect 405328 270098 405370 270334
rect 405606 270098 405648 270334
rect 405328 270014 405648 270098
rect 405328 269778 405370 270014
rect 405606 269778 405648 270014
rect 405328 269746 405648 269778
rect 338768 266614 339088 266646
rect 338768 266378 338810 266614
rect 339046 266378 339088 266614
rect 338768 266294 339088 266378
rect 338768 266058 338810 266294
rect 339046 266058 339088 266294
rect 338768 266026 339088 266058
rect 369488 266614 369808 266646
rect 369488 266378 369530 266614
rect 369766 266378 369808 266614
rect 369488 266294 369808 266378
rect 369488 266058 369530 266294
rect 369766 266058 369808 266294
rect 369488 266026 369808 266058
rect 400208 266614 400528 266646
rect 400208 266378 400250 266614
rect 400486 266378 400528 266614
rect 400208 266294 400528 266378
rect 400208 266058 400250 266294
rect 400486 266058 400528 266294
rect 400208 266026 400528 266058
rect 333648 262894 333968 262926
rect 333648 262658 333690 262894
rect 333926 262658 333968 262894
rect 333648 262574 333968 262658
rect 333648 262338 333690 262574
rect 333926 262338 333968 262574
rect 333648 262306 333968 262338
rect 364368 262894 364688 262926
rect 364368 262658 364410 262894
rect 364646 262658 364688 262894
rect 364368 262574 364688 262658
rect 364368 262338 364410 262574
rect 364646 262338 364688 262574
rect 364368 262306 364688 262338
rect 395088 262894 395408 262926
rect 395088 262658 395130 262894
rect 395366 262658 395408 262894
rect 395088 262574 395408 262658
rect 395088 262338 395130 262574
rect 395366 262338 395408 262574
rect 395088 262306 395408 262338
rect 328528 259174 328848 259206
rect 328528 258938 328570 259174
rect 328806 258938 328848 259174
rect 328528 258854 328848 258938
rect 328528 258618 328570 258854
rect 328806 258618 328848 258854
rect 328528 258586 328848 258618
rect 359248 259174 359568 259206
rect 359248 258938 359290 259174
rect 359526 258938 359568 259174
rect 359248 258854 359568 258938
rect 359248 258618 359290 258854
rect 359526 258618 359568 258854
rect 359248 258586 359568 258618
rect 389968 259174 390288 259206
rect 389968 258938 390010 259174
rect 390246 258938 390288 259174
rect 389968 258854 390288 258938
rect 389968 258618 390010 258854
rect 390246 258618 390288 258854
rect 389968 258586 390288 258618
rect 420688 259174 421008 259206
rect 420688 258938 420730 259174
rect 420966 258938 421008 259174
rect 420688 258854 421008 258938
rect 420688 258618 420730 258854
rect 420966 258618 421008 258854
rect 420688 258586 421008 258618
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 313168 234334 313488 234366
rect 313168 234098 313210 234334
rect 313446 234098 313488 234334
rect 313168 234014 313488 234098
rect 313168 233778 313210 234014
rect 313446 233778 313488 234014
rect 313168 233746 313488 233778
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 308048 194614 308368 194646
rect 308048 194378 308090 194614
rect 308326 194378 308368 194614
rect 308048 194294 308368 194378
rect 308048 194058 308090 194294
rect 308326 194058 308368 194294
rect 308048 194026 308368 194058
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 302928 154894 303248 154926
rect 302928 154658 302970 154894
rect 303206 154658 303248 154894
rect 302928 154574 303248 154658
rect 302928 154338 302970 154574
rect 303206 154338 303248 154574
rect 302928 154306 303248 154338
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 287568 94054 287888 94086
rect 287568 93818 287610 94054
rect 287846 93818 287888 94054
rect 287568 93734 287888 93818
rect 287568 93498 287610 93734
rect 287846 93498 287888 93734
rect 287568 93466 287888 93498
rect 282448 90334 282768 90366
rect 282448 90098 282490 90334
rect 282726 90098 282768 90334
rect 282448 90014 282768 90098
rect 282448 89778 282490 90014
rect 282726 89778 282768 90014
rect 282448 89746 282768 89778
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 277328 50614 277648 50646
rect 277328 50378 277370 50614
rect 277606 50378 277648 50614
rect 277328 50294 277648 50378
rect 277328 50058 277370 50294
rect 277606 50058 277648 50294
rect 277328 50026 277648 50058
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 272208 10894 272528 10926
rect 272208 10658 272250 10894
rect 272486 10658 272528 10894
rect 272208 10574 272528 10658
rect 272208 10338 272250 10574
rect 272486 10338 272528 10574
rect 272208 10306 272528 10338
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 -5146 273014 2988
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 -6106 276734 25218
rect 279834 29494 280454 64938
rect 289794 75454 290414 110898
rect 292688 111454 293008 111486
rect 292688 111218 292730 111454
rect 292966 111218 293008 111454
rect 292688 111134 293008 111218
rect 292688 110898 292730 111134
rect 292966 110898 293008 111134
rect 292688 110866 293008 110898
rect 293514 79174 294134 114618
rect 297808 115174 298128 115206
rect 297808 114938 297850 115174
rect 298086 114938 298128 115174
rect 297808 114854 298128 114938
rect 297808 114618 297850 114854
rect 298086 114618 298128 114854
rect 297808 114586 298128 114618
rect 300954 86614 301574 122058
rect 304674 126334 305294 161778
rect 312114 169774 312734 205218
rect 315834 209494 316454 244938
rect 318288 238054 318608 238086
rect 318288 237818 318330 238054
rect 318566 237818 318608 238054
rect 318288 237734 318608 237818
rect 318288 237498 318330 237734
rect 318566 237498 318608 237734
rect 318288 237466 318608 237498
rect 323408 219454 323728 219486
rect 323408 219218 323450 219454
rect 323686 219218 323728 219454
rect 323408 219134 323728 219218
rect 323408 218898 323450 219134
rect 323686 218898 323728 219134
rect 323408 218866 323728 218898
rect 325794 219454 326414 254898
rect 354128 255454 354448 255486
rect 354128 255218 354170 255454
rect 354406 255218 354448 255454
rect 354128 255134 354448 255218
rect 354128 254898 354170 255134
rect 354406 254898 354448 255134
rect 354128 254866 354448 254898
rect 384848 255454 385168 255486
rect 384848 255218 384890 255454
rect 385126 255218 385168 255454
rect 384848 255134 385168 255218
rect 384848 254898 384890 255134
rect 385126 254898 385168 255134
rect 384848 254866 385168 254898
rect 415568 255454 415888 255486
rect 415568 255218 415610 255454
rect 415846 255218 415888 255454
rect 415568 255134 415888 255218
rect 415568 254898 415610 255134
rect 415846 254898 415888 255134
rect 415568 254866 415888 254898
rect 423834 245494 424454 280938
rect 433794 291454 434414 326898
rect 437514 331174 438134 366618
rect 444954 374614 445574 410058
rect 448674 414334 449294 449778
rect 452394 454054 453014 489498
rect 459834 497494 460454 532938
rect 469794 543454 470414 578898
rect 473514 583174 474134 618618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 602500 477854 622338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 471888 562054 472208 562086
rect 471888 561818 471930 562054
rect 472166 561818 472208 562054
rect 471888 561734 472208 561818
rect 471888 561498 471930 561734
rect 472166 561498 472208 561734
rect 471888 561466 472208 561498
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 466768 522334 467088 522366
rect 466768 522098 466810 522334
rect 467046 522098 467088 522334
rect 466768 522014 467088 522098
rect 466768 521778 466810 522014
rect 467046 521778 467088 522014
rect 466768 521746 467088 521778
rect 461648 518614 461968 518646
rect 461648 518378 461690 518614
rect 461926 518378 461968 518614
rect 461648 518294 461968 518378
rect 461648 518058 461690 518294
rect 461926 518058 461968 518294
rect 461648 518026 461968 518058
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 456528 478894 456848 478926
rect 456528 478658 456570 478894
rect 456806 478658 456848 478894
rect 456528 478574 456848 478658
rect 456528 478338 456570 478574
rect 456806 478338 456848 478574
rect 456528 478306 456848 478338
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 451408 439174 451728 439206
rect 451408 438938 451450 439174
rect 451686 438938 451728 439174
rect 451408 438854 451728 438938
rect 451408 438618 451450 438854
rect 451686 438618 451728 438854
rect 451408 438586 451728 438618
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 446288 399454 446608 399486
rect 446288 399218 446330 399454
rect 446566 399218 446608 399454
rect 446288 399134 446608 399218
rect 446288 398898 446330 399134
rect 446566 398898 446608 399134
rect 446288 398866 446608 398898
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 441168 346054 441488 346086
rect 441168 345818 441210 346054
rect 441446 345818 441488 346054
rect 441168 345734 441488 345818
rect 441168 345498 441210 345734
rect 441446 345498 441488 345734
rect 441168 345466 441488 345498
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 436048 306334 436368 306366
rect 436048 306098 436090 306334
rect 436326 306098 436368 306334
rect 436048 306014 436368 306098
rect 436048 305778 436090 306014
rect 436326 305778 436368 306014
rect 436048 305746 436368 305778
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 430928 266614 431248 266646
rect 430928 266378 430970 266614
rect 431206 266378 431248 266614
rect 430928 266294 431248 266378
rect 430928 266058 430970 266294
rect 431206 266058 431248 266294
rect 430928 266026 431248 266058
rect 425808 262894 426128 262926
rect 425808 262658 425850 262894
rect 426086 262658 426128 262894
rect 425808 262574 426128 262658
rect 425808 262338 425850 262574
rect 426086 262338 426128 262574
rect 425808 262306 426128 262338
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 349008 238054 349328 238086
rect 349008 237818 349050 238054
rect 349286 237818 349328 238054
rect 349008 237734 349328 237818
rect 349008 237498 349050 237734
rect 349286 237498 349328 237734
rect 349008 237466 349328 237498
rect 379728 238054 380048 238086
rect 379728 237818 379770 238054
rect 380006 237818 380048 238054
rect 379728 237734 380048 237818
rect 379728 237498 379770 237734
rect 380006 237498 380048 237734
rect 379728 237466 380048 237498
rect 410448 238054 410768 238086
rect 410448 237818 410490 238054
rect 410726 237818 410768 238054
rect 410448 237734 410768 237818
rect 410448 237498 410490 237734
rect 410726 237498 410768 237734
rect 410448 237466 410768 237498
rect 343888 234334 344208 234366
rect 343888 234098 343930 234334
rect 344166 234098 344208 234334
rect 343888 234014 344208 234098
rect 343888 233778 343930 234014
rect 344166 233778 344208 234014
rect 343888 233746 344208 233778
rect 374608 234334 374928 234366
rect 374608 234098 374650 234334
rect 374886 234098 374928 234334
rect 374608 234014 374928 234098
rect 374608 233778 374650 234014
rect 374886 233778 374928 234014
rect 374608 233746 374928 233778
rect 405328 234334 405648 234366
rect 405328 234098 405370 234334
rect 405606 234098 405648 234334
rect 405328 234014 405648 234098
rect 405328 233778 405370 234014
rect 405606 233778 405648 234014
rect 405328 233746 405648 233778
rect 338768 230614 339088 230646
rect 338768 230378 338810 230614
rect 339046 230378 339088 230614
rect 338768 230294 339088 230378
rect 338768 230058 338810 230294
rect 339046 230058 339088 230294
rect 338768 230026 339088 230058
rect 369488 230614 369808 230646
rect 369488 230378 369530 230614
rect 369766 230378 369808 230614
rect 369488 230294 369808 230378
rect 369488 230058 369530 230294
rect 369766 230058 369808 230294
rect 369488 230026 369808 230058
rect 400208 230614 400528 230646
rect 400208 230378 400250 230614
rect 400486 230378 400528 230614
rect 400208 230294 400528 230378
rect 400208 230058 400250 230294
rect 400486 230058 400528 230294
rect 400208 230026 400528 230058
rect 333648 226894 333968 226926
rect 333648 226658 333690 226894
rect 333926 226658 333968 226894
rect 333648 226574 333968 226658
rect 333648 226338 333690 226574
rect 333926 226338 333968 226574
rect 333648 226306 333968 226338
rect 364368 226894 364688 226926
rect 364368 226658 364410 226894
rect 364646 226658 364688 226894
rect 364368 226574 364688 226658
rect 364368 226338 364410 226574
rect 364646 226338 364688 226574
rect 364368 226306 364688 226338
rect 395088 226894 395408 226926
rect 395088 226658 395130 226894
rect 395366 226658 395408 226894
rect 395088 226574 395408 226658
rect 395088 226338 395130 226574
rect 395366 226338 395408 226574
rect 395088 226306 395408 226338
rect 328528 223174 328848 223206
rect 328528 222938 328570 223174
rect 328806 222938 328848 223174
rect 328528 222854 328848 222938
rect 328528 222618 328570 222854
rect 328806 222618 328848 222854
rect 328528 222586 328848 222618
rect 359248 223174 359568 223206
rect 359248 222938 359290 223174
rect 359526 222938 359568 223174
rect 359248 222854 359568 222938
rect 359248 222618 359290 222854
rect 359526 222618 359568 222854
rect 359248 222586 359568 222618
rect 389968 223174 390288 223206
rect 389968 222938 390010 223174
rect 390246 222938 390288 223174
rect 389968 222854 390288 222938
rect 389968 222618 390010 222854
rect 390246 222618 390288 222854
rect 389968 222586 390288 222618
rect 420688 223174 421008 223206
rect 420688 222938 420730 223174
rect 420966 222938 421008 223174
rect 420688 222854 421008 222938
rect 420688 222618 420730 222854
rect 420966 222618 421008 222854
rect 420688 222586 421008 222618
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 313168 198334 313488 198366
rect 313168 198098 313210 198334
rect 313446 198098 313488 198334
rect 313168 198014 313488 198098
rect 313168 197778 313210 198014
rect 313446 197778 313488 198014
rect 313168 197746 313488 197778
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 308048 158614 308368 158646
rect 308048 158378 308090 158614
rect 308326 158378 308368 158614
rect 308048 158294 308368 158378
rect 308048 158058 308090 158294
rect 308326 158058 308368 158294
rect 308048 158026 308368 158058
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 302928 118894 303248 118926
rect 302928 118658 302970 118894
rect 303206 118658 303248 118894
rect 302928 118574 303248 118658
rect 302928 118338 302970 118574
rect 303206 118338 303248 118574
rect 302928 118306 303248 118338
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 287568 58054 287888 58086
rect 287568 57818 287610 58054
rect 287846 57818 287888 58054
rect 287568 57734 287888 57818
rect 287568 57498 287610 57734
rect 287846 57498 287888 57734
rect 287568 57466 287888 57498
rect 282448 54334 282768 54366
rect 282448 54098 282490 54334
rect 282726 54098 282768 54334
rect 282448 54014 282768 54098
rect 282448 53778 282490 54014
rect 282726 53778 282768 54014
rect 282448 53746 282768 53778
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 277328 14614 277648 14646
rect 277328 14378 277370 14614
rect 277606 14378 277648 14614
rect 277328 14294 277648 14378
rect 277328 14058 277370 14294
rect 277606 14058 277648 14294
rect 277328 14026 277648 14058
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 -7066 280454 28938
rect 289794 39454 290414 74898
rect 292688 75454 293008 75486
rect 292688 75218 292730 75454
rect 292966 75218 293008 75454
rect 292688 75134 293008 75218
rect 292688 74898 292730 75134
rect 292966 74898 293008 75134
rect 292688 74866 293008 74898
rect 293514 43174 294134 78618
rect 297808 79174 298128 79206
rect 297808 78938 297850 79174
rect 298086 78938 298128 79174
rect 297808 78854 298128 78938
rect 297808 78618 297850 78854
rect 298086 78618 298128 78854
rect 297808 78586 298128 78618
rect 300954 50614 301574 86058
rect 304674 90334 305294 125778
rect 312114 133774 312734 169218
rect 315834 173494 316454 208938
rect 318288 202054 318608 202086
rect 318288 201818 318330 202054
rect 318566 201818 318608 202054
rect 318288 201734 318608 201818
rect 318288 201498 318330 201734
rect 318566 201498 318608 201734
rect 318288 201466 318608 201498
rect 323408 183454 323728 183486
rect 323408 183218 323450 183454
rect 323686 183218 323728 183454
rect 323408 183134 323728 183218
rect 323408 182898 323450 183134
rect 323686 182898 323728 183134
rect 323408 182866 323728 182898
rect 325794 183454 326414 218898
rect 354128 219454 354448 219486
rect 354128 219218 354170 219454
rect 354406 219218 354448 219454
rect 354128 219134 354448 219218
rect 354128 218898 354170 219134
rect 354406 218898 354448 219134
rect 354128 218866 354448 218898
rect 384848 219454 385168 219486
rect 384848 219218 384890 219454
rect 385126 219218 385168 219454
rect 384848 219134 385168 219218
rect 384848 218898 384890 219134
rect 385126 218898 385168 219134
rect 384848 218866 385168 218898
rect 415568 219454 415888 219486
rect 415568 219218 415610 219454
rect 415846 219218 415888 219454
rect 415568 219134 415888 219218
rect 415568 218898 415610 219134
rect 415846 218898 415888 219134
rect 415568 218866 415888 218898
rect 423834 209494 424454 244938
rect 433794 255454 434414 290898
rect 437514 295174 438134 330618
rect 444954 338614 445574 374058
rect 448674 378334 449294 413778
rect 452394 418054 453014 453498
rect 459834 461494 460454 496938
rect 469794 507454 470414 542898
rect 473514 547174 474134 582618
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 477008 579454 477328 579486
rect 477008 579218 477050 579454
rect 477286 579218 477328 579454
rect 477008 579134 477328 579218
rect 477008 578898 477050 579134
rect 477286 578898 477328 579134
rect 477008 578866 477328 578898
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 471888 526054 472208 526086
rect 471888 525818 471930 526054
rect 472166 525818 472208 526054
rect 471888 525734 472208 525818
rect 471888 525498 471930 525734
rect 472166 525498 472208 525734
rect 471888 525466 472208 525498
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 466768 486334 467088 486366
rect 466768 486098 466810 486334
rect 467046 486098 467088 486334
rect 466768 486014 467088 486098
rect 466768 485778 466810 486014
rect 467046 485778 467088 486014
rect 466768 485746 467088 485778
rect 461648 482614 461968 482646
rect 461648 482378 461690 482614
rect 461926 482378 461968 482614
rect 461648 482294 461968 482378
rect 461648 482058 461690 482294
rect 461926 482058 461968 482294
rect 461648 482026 461968 482058
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 456528 442894 456848 442926
rect 456528 442658 456570 442894
rect 456806 442658 456848 442894
rect 456528 442574 456848 442658
rect 456528 442338 456570 442574
rect 456806 442338 456848 442574
rect 456528 442306 456848 442338
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 451408 403174 451728 403206
rect 451408 402938 451450 403174
rect 451686 402938 451728 403174
rect 451408 402854 451728 402938
rect 451408 402618 451450 402854
rect 451686 402618 451728 402854
rect 451408 402586 451728 402618
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 446288 363454 446608 363486
rect 446288 363218 446330 363454
rect 446566 363218 446608 363454
rect 446288 363134 446608 363218
rect 446288 362898 446330 363134
rect 446566 362898 446608 363134
rect 446288 362866 446608 362898
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 441168 310054 441488 310086
rect 441168 309818 441210 310054
rect 441446 309818 441488 310054
rect 441168 309734 441488 309818
rect 441168 309498 441210 309734
rect 441446 309498 441488 309734
rect 441168 309466 441488 309498
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 436048 270334 436368 270366
rect 436048 270098 436090 270334
rect 436326 270098 436368 270334
rect 436048 270014 436368 270098
rect 436048 269778 436090 270014
rect 436326 269778 436368 270014
rect 436048 269746 436368 269778
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 430928 230614 431248 230646
rect 430928 230378 430970 230614
rect 431206 230378 431248 230614
rect 430928 230294 431248 230378
rect 430928 230058 430970 230294
rect 431206 230058 431248 230294
rect 430928 230026 431248 230058
rect 425808 226894 426128 226926
rect 425808 226658 425850 226894
rect 426086 226658 426128 226894
rect 425808 226574 426128 226658
rect 425808 226338 425850 226574
rect 426086 226338 426128 226574
rect 425808 226306 426128 226338
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 349008 202054 349328 202086
rect 349008 201818 349050 202054
rect 349286 201818 349328 202054
rect 349008 201734 349328 201818
rect 349008 201498 349050 201734
rect 349286 201498 349328 201734
rect 349008 201466 349328 201498
rect 379728 202054 380048 202086
rect 379728 201818 379770 202054
rect 380006 201818 380048 202054
rect 379728 201734 380048 201818
rect 379728 201498 379770 201734
rect 380006 201498 380048 201734
rect 379728 201466 380048 201498
rect 410448 202054 410768 202086
rect 410448 201818 410490 202054
rect 410726 201818 410768 202054
rect 410448 201734 410768 201818
rect 410448 201498 410490 201734
rect 410726 201498 410768 201734
rect 410448 201466 410768 201498
rect 343888 198334 344208 198366
rect 343888 198098 343930 198334
rect 344166 198098 344208 198334
rect 343888 198014 344208 198098
rect 343888 197778 343930 198014
rect 344166 197778 344208 198014
rect 343888 197746 344208 197778
rect 374608 198334 374928 198366
rect 374608 198098 374650 198334
rect 374886 198098 374928 198334
rect 374608 198014 374928 198098
rect 374608 197778 374650 198014
rect 374886 197778 374928 198014
rect 374608 197746 374928 197778
rect 338768 194614 339088 194646
rect 338768 194378 338810 194614
rect 339046 194378 339088 194614
rect 338768 194294 339088 194378
rect 338768 194058 338810 194294
rect 339046 194058 339088 194294
rect 338768 194026 339088 194058
rect 369488 194614 369808 194646
rect 369488 194378 369530 194614
rect 369766 194378 369808 194614
rect 369488 194294 369808 194378
rect 369488 194058 369530 194294
rect 369766 194058 369808 194294
rect 369488 194026 369808 194058
rect 400208 194431 400528 194600
rect 400208 194195 400250 194431
rect 400486 194195 400528 194431
rect 400208 194026 400528 194195
rect 333648 190894 333968 190926
rect 333648 190658 333690 190894
rect 333926 190658 333968 190894
rect 333648 190574 333968 190658
rect 333648 190338 333690 190574
rect 333926 190338 333968 190574
rect 333648 190306 333968 190338
rect 364368 190894 364688 190926
rect 364368 190658 364410 190894
rect 364646 190658 364688 190894
rect 364368 190574 364688 190658
rect 364368 190338 364410 190574
rect 364646 190338 364688 190574
rect 364368 190306 364688 190338
rect 395088 190894 395408 190926
rect 395088 190658 395130 190894
rect 395366 190658 395408 190894
rect 395088 190574 395408 190658
rect 395088 190338 395130 190574
rect 395366 190338 395408 190574
rect 395088 190306 395408 190338
rect 328528 187174 328848 187206
rect 328528 186938 328570 187174
rect 328806 186938 328848 187174
rect 328528 186854 328848 186938
rect 328528 186618 328570 186854
rect 328806 186618 328848 186854
rect 328528 186586 328848 186618
rect 359248 187174 359568 187206
rect 359248 186938 359290 187174
rect 359526 186938 359568 187174
rect 359248 186854 359568 186938
rect 359248 186618 359290 186854
rect 359526 186618 359568 186854
rect 359248 186586 359568 186618
rect 389968 187174 390288 187206
rect 389968 186938 390010 187174
rect 390246 186938 390288 187174
rect 389968 186854 390288 186938
rect 389968 186618 390010 186854
rect 390246 186618 390288 186854
rect 389968 186586 390288 186618
rect 420688 187174 421008 187206
rect 420688 186938 420730 187174
rect 420966 186938 421008 187174
rect 420688 186854 421008 186938
rect 420688 186618 420730 186854
rect 420966 186618 421008 186854
rect 420688 186586 421008 186618
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 313168 162334 313488 162366
rect 313168 162098 313210 162334
rect 313446 162098 313488 162334
rect 313168 162014 313488 162098
rect 313168 161778 313210 162014
rect 313446 161778 313488 162014
rect 313168 161746 313488 161778
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 308048 122614 308368 122646
rect 308048 122378 308090 122614
rect 308326 122378 308368 122614
rect 308048 122294 308368 122378
rect 308048 122058 308090 122294
rect 308326 122058 308368 122294
rect 308048 122026 308368 122058
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 302928 82894 303248 82926
rect 302928 82658 302970 82894
rect 303206 82658 303248 82894
rect 302928 82574 303248 82658
rect 302928 82338 302970 82574
rect 303206 82338 303248 82574
rect 302928 82306 303248 82338
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 287568 22054 287888 22086
rect 287568 21818 287610 22054
rect 287846 21818 287888 22054
rect 287568 21734 287888 21818
rect 287568 21498 287610 21734
rect 287846 21498 287888 21734
rect 287568 21466 287888 21498
rect 282448 18334 282768 18366
rect 282448 18098 282490 18334
rect 282726 18098 282768 18334
rect 282448 18014 282768 18098
rect 282448 17778 282490 18014
rect 282726 17778 282768 18014
rect 282448 17746 282768 17778
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 3454 290414 38898
rect 292688 39454 293008 39486
rect 292688 39218 292730 39454
rect 292966 39218 293008 39454
rect 292688 39134 293008 39218
rect 292688 38898 292730 39134
rect 292966 38898 293008 39134
rect 292688 38866 293008 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 42618
rect 297808 43174 298128 43206
rect 297808 42938 297850 43174
rect 298086 42938 298128 43174
rect 297808 42854 298128 42938
rect 297808 42618 297850 42854
rect 298086 42618 298128 42854
rect 297808 42586 298128 42618
rect 300954 14614 301574 50058
rect 304674 54334 305294 89778
rect 312114 97774 312734 133218
rect 315834 137494 316454 172938
rect 318288 166054 318608 166086
rect 318288 165818 318330 166054
rect 318566 165818 318608 166054
rect 318288 165734 318608 165818
rect 318288 165498 318330 165734
rect 318566 165498 318608 165734
rect 318288 165466 318608 165498
rect 323408 147454 323728 147486
rect 323408 147218 323450 147454
rect 323686 147218 323728 147454
rect 323408 147134 323728 147218
rect 323408 146898 323450 147134
rect 323686 146898 323728 147134
rect 323408 146866 323728 146898
rect 325794 147454 326414 182898
rect 354128 183454 354448 183486
rect 354128 183218 354170 183454
rect 354406 183218 354448 183454
rect 354128 183134 354448 183218
rect 354128 182898 354170 183134
rect 354406 182898 354448 183134
rect 354128 182866 354448 182898
rect 384848 183454 385168 183486
rect 384848 183218 384890 183454
rect 385126 183218 385168 183454
rect 384848 183134 385168 183218
rect 384848 182898 384890 183134
rect 385126 182898 385168 183134
rect 384848 182866 385168 182898
rect 415568 183454 415888 183486
rect 415568 183218 415610 183454
rect 415846 183218 415888 183454
rect 415568 183134 415888 183218
rect 415568 182898 415610 183134
rect 415846 182898 415888 183134
rect 415568 182866 415888 182898
rect 423834 173494 424454 208938
rect 433794 219454 434414 254898
rect 437514 259174 438134 294618
rect 444954 302614 445574 338058
rect 448674 342334 449294 377778
rect 452394 382054 453014 417498
rect 459834 425494 460454 460938
rect 469794 471454 470414 506898
rect 473514 511174 474134 546618
rect 480954 554614 481574 590058
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 630334 485294 665778
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 482128 583174 482448 583206
rect 482128 582938 482170 583174
rect 482406 582938 482448 583174
rect 482128 582854 482448 582938
rect 482128 582618 482170 582854
rect 482406 582618 482448 582854
rect 482128 582586 482448 582618
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 477008 543454 477328 543486
rect 477008 543218 477050 543454
rect 477286 543218 477328 543454
rect 477008 543134 477328 543218
rect 477008 542898 477050 543134
rect 477286 542898 477328 543134
rect 477008 542866 477328 542898
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 471888 490054 472208 490086
rect 471888 489818 471930 490054
rect 472166 489818 472208 490054
rect 471888 489734 472208 489818
rect 471888 489498 471930 489734
rect 472166 489498 472208 489734
rect 471888 489466 472208 489498
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 466768 450334 467088 450366
rect 466768 450098 466810 450334
rect 467046 450098 467088 450334
rect 466768 450014 467088 450098
rect 466768 449778 466810 450014
rect 467046 449778 467088 450014
rect 466768 449746 467088 449778
rect 461648 446614 461968 446646
rect 461648 446378 461690 446614
rect 461926 446378 461968 446614
rect 461648 446294 461968 446378
rect 461648 446058 461690 446294
rect 461926 446058 461968 446294
rect 461648 446026 461968 446058
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 456528 406894 456848 406926
rect 456528 406658 456570 406894
rect 456806 406658 456848 406894
rect 456528 406574 456848 406658
rect 456528 406338 456570 406574
rect 456806 406338 456848 406574
rect 456528 406306 456848 406338
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 451408 367174 451728 367206
rect 451408 366938 451450 367174
rect 451686 366938 451728 367174
rect 451408 366854 451728 366938
rect 451408 366618 451450 366854
rect 451686 366618 451728 366854
rect 451408 366586 451728 366618
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 446288 327454 446608 327486
rect 446288 327218 446330 327454
rect 446566 327218 446608 327454
rect 446288 327134 446608 327218
rect 446288 326898 446330 327134
rect 446566 326898 446608 327134
rect 446288 326866 446608 326898
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 441168 274054 441488 274086
rect 441168 273818 441210 274054
rect 441446 273818 441488 274054
rect 441168 273734 441488 273818
rect 441168 273498 441210 273734
rect 441446 273498 441488 273734
rect 441168 273466 441488 273498
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 436048 234334 436368 234366
rect 436048 234098 436090 234334
rect 436326 234098 436368 234334
rect 436048 234014 436368 234098
rect 436048 233778 436090 234014
rect 436326 233778 436368 234014
rect 436048 233746 436368 233778
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 430928 194614 431248 194646
rect 430928 194378 430970 194614
rect 431206 194378 431248 194614
rect 430928 194294 431248 194378
rect 430928 194058 430970 194294
rect 431206 194058 431248 194294
rect 430928 194026 431248 194058
rect 425808 190894 426128 190926
rect 425808 190658 425850 190894
rect 426086 190658 426128 190894
rect 425808 190574 426128 190658
rect 425808 190338 425850 190574
rect 426086 190338 426128 190574
rect 425808 190306 426128 190338
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 349008 166054 349328 166086
rect 349008 165818 349050 166054
rect 349286 165818 349328 166054
rect 349008 165734 349328 165818
rect 349008 165498 349050 165734
rect 349286 165498 349328 165734
rect 349008 165466 349328 165498
rect 379728 166054 380048 166086
rect 379728 165818 379770 166054
rect 380006 165818 380048 166054
rect 379728 165734 380048 165818
rect 379728 165498 379770 165734
rect 380006 165498 380048 165734
rect 379728 165466 380048 165498
rect 410448 166054 410768 166086
rect 410448 165818 410490 166054
rect 410726 165818 410768 166054
rect 410448 165734 410768 165818
rect 410448 165498 410490 165734
rect 410726 165498 410768 165734
rect 410448 165466 410768 165498
rect 343888 162334 344208 162366
rect 343888 162098 343930 162334
rect 344166 162098 344208 162334
rect 343888 162014 344208 162098
rect 343888 161778 343930 162014
rect 344166 161778 344208 162014
rect 343888 161746 344208 161778
rect 374608 162334 374928 162366
rect 374608 162098 374650 162334
rect 374886 162098 374928 162334
rect 374608 162014 374928 162098
rect 374608 161778 374650 162014
rect 374886 161778 374928 162014
rect 374608 161746 374928 161778
rect 405328 162334 405648 162366
rect 405328 162098 405370 162334
rect 405606 162098 405648 162334
rect 405328 162014 405648 162098
rect 405328 161778 405370 162014
rect 405606 161778 405648 162014
rect 405328 161746 405648 161778
rect 338768 158614 339088 158646
rect 338768 158378 338810 158614
rect 339046 158378 339088 158614
rect 338768 158294 339088 158378
rect 338768 158058 338810 158294
rect 339046 158058 339088 158294
rect 338768 158026 339088 158058
rect 369488 158614 369808 158646
rect 369488 158378 369530 158614
rect 369766 158378 369808 158614
rect 369488 158294 369808 158378
rect 369488 158058 369530 158294
rect 369766 158058 369808 158294
rect 369488 158026 369808 158058
rect 400208 158614 400528 158646
rect 400208 158378 400250 158614
rect 400486 158378 400528 158614
rect 400208 158294 400528 158378
rect 400208 158058 400250 158294
rect 400486 158058 400528 158294
rect 400208 158026 400528 158058
rect 333648 154894 333968 154926
rect 333648 154658 333690 154894
rect 333926 154658 333968 154894
rect 333648 154574 333968 154658
rect 333648 154338 333690 154574
rect 333926 154338 333968 154574
rect 333648 154306 333968 154338
rect 364368 154894 364688 154926
rect 364368 154658 364410 154894
rect 364646 154658 364688 154894
rect 364368 154574 364688 154658
rect 364368 154338 364410 154574
rect 364646 154338 364688 154574
rect 364368 154306 364688 154338
rect 395088 154894 395408 154926
rect 395088 154658 395130 154894
rect 395366 154658 395408 154894
rect 395088 154574 395408 154658
rect 395088 154338 395130 154574
rect 395366 154338 395408 154574
rect 395088 154306 395408 154338
rect 328528 151174 328848 151206
rect 328528 150938 328570 151174
rect 328806 150938 328848 151174
rect 328528 150854 328848 150938
rect 328528 150618 328570 150854
rect 328806 150618 328848 150854
rect 328528 150586 328848 150618
rect 359248 151174 359568 151206
rect 359248 150938 359290 151174
rect 359526 150938 359568 151174
rect 359248 150854 359568 150938
rect 359248 150618 359290 150854
rect 359526 150618 359568 150854
rect 359248 150586 359568 150618
rect 389968 151174 390288 151206
rect 389968 150938 390010 151174
rect 390246 150938 390288 151174
rect 389968 150854 390288 150938
rect 389968 150618 390010 150854
rect 390246 150618 390288 150854
rect 389968 150586 390288 150618
rect 420688 151174 421008 151206
rect 420688 150938 420730 151174
rect 420966 150938 421008 151174
rect 420688 150854 421008 150938
rect 420688 150618 420730 150854
rect 420966 150618 421008 150854
rect 420688 150586 421008 150618
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 313168 126334 313488 126366
rect 313168 126098 313210 126334
rect 313446 126098 313488 126334
rect 313168 126014 313488 126098
rect 313168 125778 313210 126014
rect 313446 125778 313488 126014
rect 313168 125746 313488 125778
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 308048 86614 308368 86646
rect 308048 86378 308090 86614
rect 308326 86378 308368 86614
rect 308048 86294 308368 86378
rect 308048 86058 308090 86294
rect 308326 86058 308368 86294
rect 308048 86026 308368 86058
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 302928 46894 303248 46926
rect 302928 46658 302970 46894
rect 303206 46658 303248 46894
rect 302928 46574 303248 46658
rect 302928 46338 302970 46574
rect 303206 46338 303248 46574
rect 302928 46306 303248 46338
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 297808 7174 298128 7206
rect 297808 6938 297850 7174
rect 298086 6938 298128 7174
rect 297808 6854 298128 6938
rect 297808 6618 297850 6854
rect 298086 6618 298128 6854
rect 297808 6586 298128 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 -2266 297854 2988
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 -3226 301574 14058
rect 304674 18334 305294 53778
rect 312114 61774 312734 97218
rect 315834 101494 316454 136938
rect 318288 130054 318608 130086
rect 318288 129818 318330 130054
rect 318566 129818 318608 130054
rect 318288 129734 318608 129818
rect 318288 129498 318330 129734
rect 318566 129498 318608 129734
rect 318288 129466 318608 129498
rect 323408 111454 323728 111486
rect 323408 111218 323450 111454
rect 323686 111218 323728 111454
rect 323408 111134 323728 111218
rect 323408 110898 323450 111134
rect 323686 110898 323728 111134
rect 323408 110866 323728 110898
rect 325794 111454 326414 146898
rect 354128 147454 354448 147486
rect 354128 147218 354170 147454
rect 354406 147218 354448 147454
rect 354128 147134 354448 147218
rect 354128 146898 354170 147134
rect 354406 146898 354448 147134
rect 354128 146866 354448 146898
rect 384848 147454 385168 147486
rect 384848 147218 384890 147454
rect 385126 147218 385168 147454
rect 384848 147134 385168 147218
rect 384848 146898 384890 147134
rect 385126 146898 385168 147134
rect 384848 146866 385168 146898
rect 415568 147454 415888 147486
rect 415568 147218 415610 147454
rect 415846 147218 415888 147454
rect 415568 147134 415888 147218
rect 415568 146898 415610 147134
rect 415846 146898 415888 147134
rect 415568 146866 415888 146898
rect 423834 137494 424454 172938
rect 433794 183454 434414 218898
rect 437514 223174 438134 258618
rect 444954 266614 445574 302058
rect 448674 306334 449294 341778
rect 452394 346054 453014 381498
rect 459834 389494 460454 424938
rect 469794 435454 470414 470898
rect 473514 475174 474134 510618
rect 480954 518614 481574 554058
rect 484674 558334 485294 593778
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 634054 489014 669498
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 637774 492734 673218
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 602500 492734 637218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 641494 496454 676938
rect 495834 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 496454 641494
rect 495834 641174 496454 641258
rect 495834 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 496454 641174
rect 495834 605494 496454 640938
rect 495834 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 496454 605494
rect 495834 605174 496454 605258
rect 495834 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 496454 605174
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 487248 586894 487568 586926
rect 487248 586658 487290 586894
rect 487526 586658 487568 586894
rect 487248 586574 487568 586658
rect 487248 586338 487290 586574
rect 487526 586338 487568 586574
rect 487248 586306 487568 586338
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 482128 547174 482448 547206
rect 482128 546938 482170 547174
rect 482406 546938 482448 547174
rect 482128 546854 482448 546938
rect 482128 546618 482170 546854
rect 482406 546618 482448 546854
rect 482128 546586 482448 546618
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 477008 507454 477328 507486
rect 477008 507218 477050 507454
rect 477286 507218 477328 507454
rect 477008 507134 477328 507218
rect 477008 506898 477050 507134
rect 477286 506898 477328 507134
rect 477008 506866 477328 506898
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 471888 454054 472208 454086
rect 471888 453818 471930 454054
rect 472166 453818 472208 454054
rect 471888 453734 472208 453818
rect 471888 453498 471930 453734
rect 472166 453498 472208 453734
rect 471888 453466 472208 453498
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 466768 414334 467088 414366
rect 466768 414098 466810 414334
rect 467046 414098 467088 414334
rect 466768 414014 467088 414098
rect 466768 413778 466810 414014
rect 467046 413778 467088 414014
rect 466768 413746 467088 413778
rect 461648 410614 461968 410646
rect 461648 410378 461690 410614
rect 461926 410378 461968 410614
rect 461648 410294 461968 410378
rect 461648 410058 461690 410294
rect 461926 410058 461968 410294
rect 461648 410026 461968 410058
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 456528 370894 456848 370926
rect 456528 370658 456570 370894
rect 456806 370658 456848 370894
rect 456528 370574 456848 370658
rect 456528 370338 456570 370574
rect 456806 370338 456848 370574
rect 456528 370306 456848 370338
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 451408 331174 451728 331206
rect 451408 330938 451450 331174
rect 451686 330938 451728 331174
rect 451408 330854 451728 330938
rect 451408 330618 451450 330854
rect 451686 330618 451728 330854
rect 451408 330586 451728 330618
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 446288 291454 446608 291486
rect 446288 291218 446330 291454
rect 446566 291218 446608 291454
rect 446288 291134 446608 291218
rect 446288 290898 446330 291134
rect 446566 290898 446608 291134
rect 446288 290866 446608 290898
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 441168 238054 441488 238086
rect 441168 237818 441210 238054
rect 441446 237818 441488 238054
rect 441168 237734 441488 237818
rect 441168 237498 441210 237734
rect 441446 237498 441488 237734
rect 441168 237466 441488 237498
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 436048 198334 436368 198366
rect 436048 198098 436090 198334
rect 436326 198098 436368 198334
rect 436048 198014 436368 198098
rect 436048 197778 436090 198014
rect 436326 197778 436368 198014
rect 436048 197746 436368 197778
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 430928 158614 431248 158646
rect 430928 158378 430970 158614
rect 431206 158378 431248 158614
rect 430928 158294 431248 158378
rect 430928 158058 430970 158294
rect 431206 158058 431248 158294
rect 430928 158026 431248 158058
rect 425808 154894 426128 154926
rect 425808 154658 425850 154894
rect 426086 154658 426128 154894
rect 425808 154574 426128 154658
rect 425808 154338 425850 154574
rect 426086 154338 426128 154574
rect 425808 154306 426128 154338
rect 423834 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 424454 137494
rect 423834 137174 424454 137258
rect 423834 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 424454 137174
rect 349008 130054 349328 130086
rect 349008 129818 349050 130054
rect 349286 129818 349328 130054
rect 349008 129734 349328 129818
rect 349008 129498 349050 129734
rect 349286 129498 349328 129734
rect 349008 129466 349328 129498
rect 379728 130054 380048 130086
rect 379728 129818 379770 130054
rect 380006 129818 380048 130054
rect 379728 129734 380048 129818
rect 379728 129498 379770 129734
rect 380006 129498 380048 129734
rect 379728 129466 380048 129498
rect 410448 130054 410768 130086
rect 410448 129818 410490 130054
rect 410726 129818 410768 130054
rect 410448 129734 410768 129818
rect 410448 129498 410490 129734
rect 410726 129498 410768 129734
rect 410448 129466 410768 129498
rect 343888 126334 344208 126366
rect 343888 126098 343930 126334
rect 344166 126098 344208 126334
rect 343888 126014 344208 126098
rect 343888 125778 343930 126014
rect 344166 125778 344208 126014
rect 343888 125746 344208 125778
rect 374608 126334 374928 126366
rect 374608 126098 374650 126334
rect 374886 126098 374928 126334
rect 374608 126014 374928 126098
rect 374608 125778 374650 126014
rect 374886 125778 374928 126014
rect 374608 125746 374928 125778
rect 405328 126334 405648 126366
rect 405328 126098 405370 126334
rect 405606 126098 405648 126334
rect 405328 126014 405648 126098
rect 405328 125778 405370 126014
rect 405606 125778 405648 126014
rect 405328 125746 405648 125778
rect 338768 122614 339088 122646
rect 338768 122378 338810 122614
rect 339046 122378 339088 122614
rect 338768 122294 339088 122378
rect 338768 122058 338810 122294
rect 339046 122058 339088 122294
rect 338768 122026 339088 122058
rect 369488 122614 369808 122646
rect 369488 122378 369530 122614
rect 369766 122378 369808 122614
rect 369488 122294 369808 122378
rect 369488 122058 369530 122294
rect 369766 122058 369808 122294
rect 369488 122026 369808 122058
rect 400208 122614 400528 122646
rect 400208 122378 400250 122614
rect 400486 122378 400528 122614
rect 400208 122294 400528 122378
rect 400208 122058 400250 122294
rect 400486 122058 400528 122294
rect 400208 122026 400528 122058
rect 333648 118894 333968 118926
rect 333648 118658 333690 118894
rect 333926 118658 333968 118894
rect 333648 118574 333968 118658
rect 333648 118338 333690 118574
rect 333926 118338 333968 118574
rect 333648 118306 333968 118338
rect 364368 118894 364688 118926
rect 364368 118658 364410 118894
rect 364646 118658 364688 118894
rect 364368 118574 364688 118658
rect 364368 118338 364410 118574
rect 364646 118338 364688 118574
rect 364368 118306 364688 118338
rect 395088 118894 395408 118926
rect 395088 118658 395130 118894
rect 395366 118658 395408 118894
rect 395088 118574 395408 118658
rect 395088 118338 395130 118574
rect 395366 118338 395408 118574
rect 395088 118306 395408 118338
rect 328528 115174 328848 115206
rect 328528 114938 328570 115174
rect 328806 114938 328848 115174
rect 328528 114854 328848 114938
rect 328528 114618 328570 114854
rect 328806 114618 328848 114854
rect 328528 114586 328848 114618
rect 359248 115174 359568 115206
rect 359248 114938 359290 115174
rect 359526 114938 359568 115174
rect 359248 114854 359568 114938
rect 359248 114618 359290 114854
rect 359526 114618 359568 114854
rect 359248 114586 359568 114618
rect 389968 115174 390288 115206
rect 389968 114938 390010 115174
rect 390246 114938 390288 115174
rect 389968 114854 390288 114938
rect 389968 114618 390010 114854
rect 390246 114618 390288 114854
rect 389968 114586 390288 114618
rect 420688 115174 421008 115206
rect 420688 114938 420730 115174
rect 420966 114938 421008 115174
rect 420688 114854 421008 114938
rect 420688 114618 420730 114854
rect 420966 114618 421008 114854
rect 420688 114586 421008 114618
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 313168 90334 313488 90366
rect 313168 90098 313210 90334
rect 313446 90098 313488 90334
rect 313168 90014 313488 90098
rect 313168 89778 313210 90014
rect 313446 89778 313488 90014
rect 313168 89746 313488 89778
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 308048 50614 308368 50646
rect 308048 50378 308090 50614
rect 308326 50378 308368 50614
rect 308048 50294 308368 50378
rect 308048 50058 308090 50294
rect 308326 50058 308368 50294
rect 308048 50026 308368 50058
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 302928 10894 303248 10926
rect 302928 10658 302970 10894
rect 303206 10658 303248 10894
rect 302928 10574 303248 10658
rect 302928 10338 302970 10574
rect 303206 10338 303248 10574
rect 302928 10306 303248 10338
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 -4186 305294 17778
rect 312114 25774 312734 61218
rect 315834 65494 316454 100938
rect 318288 94054 318608 94086
rect 318288 93818 318330 94054
rect 318566 93818 318608 94054
rect 318288 93734 318608 93818
rect 318288 93498 318330 93734
rect 318566 93498 318608 93734
rect 318288 93466 318608 93498
rect 323408 75454 323728 75486
rect 323408 75218 323450 75454
rect 323686 75218 323728 75454
rect 323408 75134 323728 75218
rect 323408 74898 323450 75134
rect 323686 74898 323728 75134
rect 323408 74866 323728 74898
rect 325794 75454 326414 110898
rect 354128 111454 354448 111486
rect 354128 111218 354170 111454
rect 354406 111218 354448 111454
rect 354128 111134 354448 111218
rect 354128 110898 354170 111134
rect 354406 110898 354448 111134
rect 354128 110866 354448 110898
rect 384848 111454 385168 111486
rect 384848 111218 384890 111454
rect 385126 111218 385168 111454
rect 384848 111134 385168 111218
rect 384848 110898 384890 111134
rect 385126 110898 385168 111134
rect 384848 110866 385168 110898
rect 415568 111454 415888 111486
rect 415568 111218 415610 111454
rect 415846 111218 415888 111454
rect 415568 111134 415888 111218
rect 415568 110898 415610 111134
rect 415846 110898 415888 111134
rect 415568 110866 415888 110898
rect 423834 101494 424454 136938
rect 433794 147454 434414 182898
rect 437514 187174 438134 222618
rect 444954 230614 445574 266058
rect 448674 270334 449294 305778
rect 452394 310054 453014 345498
rect 459834 353494 460454 388938
rect 469794 399454 470414 434898
rect 473514 439174 474134 474618
rect 480954 482614 481574 518058
rect 484674 522334 485294 557778
rect 488394 562054 489014 597498
rect 492368 590614 492688 590646
rect 492368 590378 492410 590614
rect 492646 590378 492688 590614
rect 492368 590294 492688 590378
rect 492368 590058 492410 590294
rect 492646 590058 492688 590294
rect 492368 590026 492688 590058
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 487248 550894 487568 550926
rect 487248 550658 487290 550894
rect 487526 550658 487568 550894
rect 487248 550574 487568 550658
rect 487248 550338 487290 550574
rect 487526 550338 487568 550574
rect 487248 550306 487568 550338
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 482128 511174 482448 511206
rect 482128 510938 482170 511174
rect 482406 510938 482448 511174
rect 482128 510854 482448 510938
rect 482128 510618 482170 510854
rect 482406 510618 482448 510854
rect 482128 510586 482448 510618
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 477008 471454 477328 471486
rect 477008 471218 477050 471454
rect 477286 471218 477328 471454
rect 477008 471134 477328 471218
rect 477008 470898 477050 471134
rect 477286 470898 477328 471134
rect 477008 470866 477328 470898
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 471888 418054 472208 418086
rect 471888 417818 471930 418054
rect 472166 417818 472208 418054
rect 471888 417734 472208 417818
rect 471888 417498 471930 417734
rect 472166 417498 472208 417734
rect 471888 417466 472208 417498
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 466768 378334 467088 378366
rect 466768 378098 466810 378334
rect 467046 378098 467088 378334
rect 466768 378014 467088 378098
rect 466768 377778 466810 378014
rect 467046 377778 467088 378014
rect 466768 377746 467088 377778
rect 461648 374614 461968 374646
rect 461648 374378 461690 374614
rect 461926 374378 461968 374614
rect 461648 374294 461968 374378
rect 461648 374058 461690 374294
rect 461926 374058 461968 374294
rect 461648 374026 461968 374058
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 456528 334894 456848 334926
rect 456528 334658 456570 334894
rect 456806 334658 456848 334894
rect 456528 334574 456848 334658
rect 456528 334338 456570 334574
rect 456806 334338 456848 334574
rect 456528 334306 456848 334338
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 451408 295174 451728 295206
rect 451408 294938 451450 295174
rect 451686 294938 451728 295174
rect 451408 294854 451728 294938
rect 451408 294618 451450 294854
rect 451686 294618 451728 294854
rect 451408 294586 451728 294618
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 446288 255454 446608 255486
rect 446288 255218 446330 255454
rect 446566 255218 446608 255454
rect 446288 255134 446608 255218
rect 446288 254898 446330 255134
rect 446566 254898 446608 255134
rect 446288 254866 446608 254898
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 441168 202054 441488 202086
rect 441168 201818 441210 202054
rect 441446 201818 441488 202054
rect 441168 201734 441488 201818
rect 441168 201498 441210 201734
rect 441446 201498 441488 201734
rect 441168 201466 441488 201498
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 436048 162334 436368 162366
rect 436048 162098 436090 162334
rect 436326 162098 436368 162334
rect 436048 162014 436368 162098
rect 436048 161778 436090 162014
rect 436326 161778 436368 162014
rect 436048 161746 436368 161778
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 430928 122614 431248 122646
rect 430928 122378 430970 122614
rect 431206 122378 431248 122614
rect 430928 122294 431248 122378
rect 430928 122058 430970 122294
rect 431206 122058 431248 122294
rect 430928 122026 431248 122058
rect 425808 118894 426128 118926
rect 425808 118658 425850 118894
rect 426086 118658 426128 118894
rect 425808 118574 426128 118658
rect 425808 118338 425850 118574
rect 426086 118338 426128 118574
rect 425808 118306 426128 118338
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 349008 94054 349328 94086
rect 349008 93818 349050 94054
rect 349286 93818 349328 94054
rect 349008 93734 349328 93818
rect 349008 93498 349050 93734
rect 349286 93498 349328 93734
rect 349008 93466 349328 93498
rect 379728 94054 380048 94086
rect 379728 93818 379770 94054
rect 380006 93818 380048 94054
rect 379728 93734 380048 93818
rect 379728 93498 379770 93734
rect 380006 93498 380048 93734
rect 379728 93466 380048 93498
rect 410448 94054 410768 94086
rect 410448 93818 410490 94054
rect 410726 93818 410768 94054
rect 410448 93734 410768 93818
rect 410448 93498 410490 93734
rect 410726 93498 410768 93734
rect 410448 93466 410768 93498
rect 343888 90334 344208 90366
rect 343888 90098 343930 90334
rect 344166 90098 344208 90334
rect 343888 90014 344208 90098
rect 343888 89778 343930 90014
rect 344166 89778 344208 90014
rect 343888 89746 344208 89778
rect 374608 90334 374928 90366
rect 374608 90098 374650 90334
rect 374886 90098 374928 90334
rect 374608 90014 374928 90098
rect 374608 89778 374650 90014
rect 374886 89778 374928 90014
rect 374608 89746 374928 89778
rect 405328 90334 405648 90366
rect 405328 90098 405370 90334
rect 405606 90098 405648 90334
rect 405328 90014 405648 90098
rect 405328 89778 405370 90014
rect 405606 89778 405648 90014
rect 405328 89746 405648 89778
rect 338768 86614 339088 86646
rect 338768 86378 338810 86614
rect 339046 86378 339088 86614
rect 338768 86294 339088 86378
rect 338768 86058 338810 86294
rect 339046 86058 339088 86294
rect 338768 86026 339088 86058
rect 369488 86614 369808 86646
rect 369488 86378 369530 86614
rect 369766 86378 369808 86614
rect 369488 86294 369808 86378
rect 369488 86058 369530 86294
rect 369766 86058 369808 86294
rect 369488 86026 369808 86058
rect 400208 86614 400528 86646
rect 400208 86378 400250 86614
rect 400486 86378 400528 86614
rect 400208 86294 400528 86378
rect 400208 86058 400250 86294
rect 400486 86058 400528 86294
rect 400208 86026 400528 86058
rect 333648 82894 333968 82926
rect 333648 82658 333690 82894
rect 333926 82658 333968 82894
rect 333648 82574 333968 82658
rect 333648 82338 333690 82574
rect 333926 82338 333968 82574
rect 333648 82306 333968 82338
rect 364368 82894 364688 82926
rect 364368 82658 364410 82894
rect 364646 82658 364688 82894
rect 364368 82574 364688 82658
rect 364368 82338 364410 82574
rect 364646 82338 364688 82574
rect 364368 82306 364688 82338
rect 395088 82894 395408 82926
rect 395088 82658 395130 82894
rect 395366 82658 395408 82894
rect 395088 82574 395408 82658
rect 395088 82338 395130 82574
rect 395366 82338 395408 82574
rect 395088 82306 395408 82338
rect 328528 79174 328848 79206
rect 328528 78938 328570 79174
rect 328806 78938 328848 79174
rect 328528 78854 328848 78938
rect 328528 78618 328570 78854
rect 328806 78618 328848 78854
rect 328528 78586 328848 78618
rect 359248 79174 359568 79206
rect 359248 78938 359290 79174
rect 359526 78938 359568 79174
rect 359248 78854 359568 78938
rect 359248 78618 359290 78854
rect 359526 78618 359568 78854
rect 359248 78586 359568 78618
rect 389968 79174 390288 79206
rect 389968 78938 390010 79174
rect 390246 78938 390288 79174
rect 389968 78854 390288 78938
rect 389968 78618 390010 78854
rect 390246 78618 390288 78854
rect 389968 78586 390288 78618
rect 420688 79174 421008 79206
rect 420688 78938 420730 79174
rect 420966 78938 421008 79174
rect 420688 78854 421008 78938
rect 420688 78618 420730 78854
rect 420966 78618 421008 78854
rect 420688 78586 421008 78618
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 313168 54334 313488 54366
rect 313168 54098 313210 54334
rect 313446 54098 313488 54334
rect 313168 54014 313488 54098
rect 313168 53778 313210 54014
rect 313446 53778 313488 54014
rect 313168 53746 313488 53778
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 308048 14614 308368 14646
rect 308048 14378 308090 14614
rect 308326 14378 308368 14614
rect 308048 14294 308368 14378
rect 308048 14058 308090 14294
rect 308326 14058 308368 14294
rect 308048 14026 308368 14058
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 -5146 309014 2988
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 -6106 312734 25218
rect 315834 29494 316454 64938
rect 318288 58054 318608 58086
rect 318288 57818 318330 58054
rect 318566 57818 318608 58054
rect 318288 57734 318608 57818
rect 318288 57498 318330 57734
rect 318566 57498 318608 57734
rect 318288 57466 318608 57498
rect 323408 39454 323728 39486
rect 323408 39218 323450 39454
rect 323686 39218 323728 39454
rect 323408 39134 323728 39218
rect 323408 38898 323450 39134
rect 323686 38898 323728 39134
rect 323408 38866 323728 38898
rect 325794 39454 326414 74898
rect 354128 75454 354448 75486
rect 354128 75218 354170 75454
rect 354406 75218 354448 75454
rect 354128 75134 354448 75218
rect 354128 74898 354170 75134
rect 354406 74898 354448 75134
rect 354128 74866 354448 74898
rect 384848 75454 385168 75486
rect 384848 75218 384890 75454
rect 385126 75218 385168 75454
rect 384848 75134 385168 75218
rect 384848 74898 384890 75134
rect 385126 74898 385168 75134
rect 384848 74866 385168 74898
rect 415568 75454 415888 75486
rect 415568 75218 415610 75454
rect 415846 75218 415888 75454
rect 415568 75134 415888 75218
rect 415568 74898 415610 75134
rect 415846 74898 415888 75134
rect 415568 74866 415888 74898
rect 423834 65494 424454 100938
rect 433794 111454 434414 146898
rect 437514 151174 438134 186618
rect 444954 194614 445574 230058
rect 448674 234334 449294 269778
rect 452394 274054 453014 309498
rect 459834 317494 460454 352938
rect 469794 363454 470414 398898
rect 473514 403174 474134 438618
rect 480954 446614 481574 482058
rect 484674 486334 485294 521778
rect 488394 526054 489014 561498
rect 495834 569494 496454 604938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 502608 598054 502928 598086
rect 502608 597818 502650 598054
rect 502886 597818 502928 598054
rect 502608 597734 502928 597818
rect 502608 597498 502650 597734
rect 502886 597498 502928 597734
rect 502608 597466 502928 597498
rect 497488 594334 497808 594366
rect 497488 594098 497530 594334
rect 497766 594098 497808 594334
rect 497488 594014 497808 594098
rect 497488 593778 497530 594014
rect 497766 593778 497808 594014
rect 497488 593746 497808 593778
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 492368 554614 492688 554646
rect 492368 554378 492410 554614
rect 492646 554378 492688 554614
rect 492368 554294 492688 554378
rect 492368 554058 492410 554294
rect 492646 554058 492688 554294
rect 492368 554026 492688 554058
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 487248 514894 487568 514926
rect 487248 514658 487290 514894
rect 487526 514658 487568 514894
rect 487248 514574 487568 514658
rect 487248 514338 487290 514574
rect 487526 514338 487568 514574
rect 487248 514306 487568 514338
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 482128 475174 482448 475206
rect 482128 474938 482170 475174
rect 482406 474938 482448 475174
rect 482128 474854 482448 474938
rect 482128 474618 482170 474854
rect 482406 474618 482448 474854
rect 482128 474586 482448 474618
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 477008 435454 477328 435486
rect 477008 435218 477050 435454
rect 477286 435218 477328 435454
rect 477008 435134 477328 435218
rect 477008 434898 477050 435134
rect 477286 434898 477328 435134
rect 477008 434866 477328 434898
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 471888 382054 472208 382086
rect 471888 381818 471930 382054
rect 472166 381818 472208 382054
rect 471888 381734 472208 381818
rect 471888 381498 471930 381734
rect 472166 381498 472208 381734
rect 471888 381466 472208 381498
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 466768 342334 467088 342366
rect 466768 342098 466810 342334
rect 467046 342098 467088 342334
rect 466768 342014 467088 342098
rect 466768 341778 466810 342014
rect 467046 341778 467088 342014
rect 466768 341746 467088 341778
rect 461648 338614 461968 338646
rect 461648 338378 461690 338614
rect 461926 338378 461968 338614
rect 461648 338294 461968 338378
rect 461648 338058 461690 338294
rect 461926 338058 461968 338294
rect 461648 338026 461968 338058
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 456528 298894 456848 298926
rect 456528 298658 456570 298894
rect 456806 298658 456848 298894
rect 456528 298574 456848 298658
rect 456528 298338 456570 298574
rect 456806 298338 456848 298574
rect 456528 298306 456848 298338
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 451408 259174 451728 259206
rect 451408 258938 451450 259174
rect 451686 258938 451728 259174
rect 451408 258854 451728 258938
rect 451408 258618 451450 258854
rect 451686 258618 451728 258854
rect 451408 258586 451728 258618
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 446288 219454 446608 219486
rect 446288 219218 446330 219454
rect 446566 219218 446608 219454
rect 446288 219134 446608 219218
rect 446288 218898 446330 219134
rect 446566 218898 446608 219134
rect 446288 218866 446608 218898
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 441168 166054 441488 166086
rect 441168 165818 441210 166054
rect 441446 165818 441488 166054
rect 441168 165734 441488 165818
rect 441168 165498 441210 165734
rect 441446 165498 441488 165734
rect 441168 165466 441488 165498
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 436048 126334 436368 126366
rect 436048 126098 436090 126334
rect 436326 126098 436368 126334
rect 436048 126014 436368 126098
rect 436048 125778 436090 126014
rect 436326 125778 436368 126014
rect 436048 125746 436368 125778
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 430928 86614 431248 86646
rect 430928 86378 430970 86614
rect 431206 86378 431248 86614
rect 430928 86294 431248 86378
rect 430928 86058 430970 86294
rect 431206 86058 431248 86294
rect 430928 86026 431248 86058
rect 425808 82894 426128 82926
rect 425808 82658 425850 82894
rect 426086 82658 426128 82894
rect 425808 82574 426128 82658
rect 425808 82338 425850 82574
rect 426086 82338 426128 82574
rect 425808 82306 426128 82338
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 349008 58054 349328 58086
rect 349008 57818 349050 58054
rect 349286 57818 349328 58054
rect 349008 57734 349328 57818
rect 349008 57498 349050 57734
rect 349286 57498 349328 57734
rect 349008 57466 349328 57498
rect 379728 58054 380048 58086
rect 379728 57818 379770 58054
rect 380006 57818 380048 58054
rect 379728 57734 380048 57818
rect 379728 57498 379770 57734
rect 380006 57498 380048 57734
rect 379728 57466 380048 57498
rect 410448 58054 410768 58086
rect 410448 57818 410490 58054
rect 410726 57818 410768 58054
rect 410448 57734 410768 57818
rect 410448 57498 410490 57734
rect 410726 57498 410768 57734
rect 410448 57466 410768 57498
rect 343888 54334 344208 54366
rect 343888 54098 343930 54334
rect 344166 54098 344208 54334
rect 343888 54014 344208 54098
rect 343888 53778 343930 54014
rect 344166 53778 344208 54014
rect 343888 53746 344208 53778
rect 374608 54334 374928 54366
rect 374608 54098 374650 54334
rect 374886 54098 374928 54334
rect 374608 54014 374928 54098
rect 374608 53778 374650 54014
rect 374886 53778 374928 54014
rect 374608 53746 374928 53778
rect 405328 54334 405648 54366
rect 405328 54098 405370 54334
rect 405606 54098 405648 54334
rect 405328 54014 405648 54098
rect 405328 53778 405370 54014
rect 405606 53778 405648 54014
rect 405328 53746 405648 53778
rect 338768 50614 339088 50646
rect 338768 50378 338810 50614
rect 339046 50378 339088 50614
rect 338768 50294 339088 50378
rect 338768 50058 338810 50294
rect 339046 50058 339088 50294
rect 338768 50026 339088 50058
rect 369488 50614 369808 50646
rect 369488 50378 369530 50614
rect 369766 50378 369808 50614
rect 369488 50294 369808 50378
rect 369488 50058 369530 50294
rect 369766 50058 369808 50294
rect 369488 50026 369808 50058
rect 400208 50614 400528 50646
rect 400208 50378 400250 50614
rect 400486 50378 400528 50614
rect 400208 50294 400528 50378
rect 400208 50058 400250 50294
rect 400486 50058 400528 50294
rect 400208 50026 400528 50058
rect 333648 46894 333968 46926
rect 333648 46658 333690 46894
rect 333926 46658 333968 46894
rect 333648 46574 333968 46658
rect 333648 46338 333690 46574
rect 333926 46338 333968 46574
rect 333648 46306 333968 46338
rect 364368 46894 364688 46926
rect 364368 46658 364410 46894
rect 364646 46658 364688 46894
rect 364368 46574 364688 46658
rect 364368 46338 364410 46574
rect 364646 46338 364688 46574
rect 364368 46306 364688 46338
rect 395088 46894 395408 46926
rect 395088 46658 395130 46894
rect 395366 46658 395408 46894
rect 395088 46574 395408 46658
rect 395088 46338 395130 46574
rect 395366 46338 395408 46574
rect 395088 46306 395408 46338
rect 328528 43174 328848 43206
rect 328528 42938 328570 43174
rect 328806 42938 328848 43174
rect 328528 42854 328848 42938
rect 328528 42618 328570 42854
rect 328806 42618 328848 42854
rect 328528 42586 328848 42618
rect 359248 43174 359568 43206
rect 359248 42938 359290 43174
rect 359526 42938 359568 43174
rect 359248 42854 359568 42938
rect 359248 42618 359290 42854
rect 359526 42618 359568 42854
rect 359248 42586 359568 42618
rect 389968 43174 390288 43206
rect 389968 42938 390010 43174
rect 390246 42938 390288 43174
rect 389968 42854 390288 42938
rect 389968 42618 390010 42854
rect 390246 42618 390288 42854
rect 389968 42586 390288 42618
rect 420688 43174 421008 43206
rect 420688 42938 420730 43174
rect 420966 42938 421008 43174
rect 420688 42854 421008 42938
rect 420688 42618 420730 42854
rect 420966 42618 421008 42854
rect 420688 42586 421008 42618
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 313168 18334 313488 18366
rect 313168 18098 313210 18334
rect 313446 18098 313488 18334
rect 313168 18014 313488 18098
rect 313168 17778 313210 18014
rect 313446 17778 313488 18014
rect 313168 17746 313488 17778
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 -7066 316454 28938
rect 318288 22054 318608 22086
rect 318288 21818 318330 22054
rect 318566 21818 318608 22054
rect 318288 21734 318608 21818
rect 318288 21498 318330 21734
rect 318566 21498 318608 21734
rect 318288 21466 318608 21498
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 3454 326414 38898
rect 354128 39454 354448 39486
rect 354128 39218 354170 39454
rect 354406 39218 354448 39454
rect 354128 39134 354448 39218
rect 354128 38898 354170 39134
rect 354406 38898 354448 39134
rect 354128 38866 354448 38898
rect 384848 39454 385168 39486
rect 384848 39218 384890 39454
rect 385126 39218 385168 39454
rect 384848 39134 385168 39218
rect 384848 38898 384890 39134
rect 385126 38898 385168 39134
rect 384848 38866 385168 38898
rect 415568 39454 415888 39486
rect 415568 39218 415610 39454
rect 415846 39218 415888 39454
rect 415568 39134 415888 39218
rect 415568 38898 415610 39134
rect 415846 38898 415888 39134
rect 415568 38866 415888 38898
rect 423834 29494 424454 64938
rect 433794 75454 434414 110898
rect 437514 115174 438134 150618
rect 444954 158614 445574 194058
rect 448674 198334 449294 233778
rect 452394 238054 453014 273498
rect 459834 281494 460454 316938
rect 469794 327454 470414 362898
rect 473514 367174 474134 402618
rect 480954 410614 481574 446058
rect 484674 450334 485294 485778
rect 488394 490054 489014 525498
rect 495834 533494 496454 568938
rect 505794 579454 506414 614898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 502608 562054 502928 562086
rect 502608 561818 502650 562054
rect 502886 561818 502928 562054
rect 502608 561734 502928 561818
rect 502608 561498 502650 561734
rect 502886 561498 502928 561734
rect 502608 561466 502928 561498
rect 497488 558334 497808 558366
rect 497488 558098 497530 558334
rect 497766 558098 497808 558334
rect 497488 558014 497808 558098
rect 497488 557778 497530 558014
rect 497766 557778 497808 558014
rect 497488 557746 497808 557778
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 492368 518614 492688 518646
rect 492368 518378 492410 518614
rect 492646 518378 492688 518614
rect 492368 518294 492688 518378
rect 492368 518058 492410 518294
rect 492646 518058 492688 518294
rect 492368 518026 492688 518058
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 487248 478894 487568 478926
rect 487248 478658 487290 478894
rect 487526 478658 487568 478894
rect 487248 478574 487568 478658
rect 487248 478338 487290 478574
rect 487526 478338 487568 478574
rect 487248 478306 487568 478338
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 482128 439174 482448 439206
rect 482128 438938 482170 439174
rect 482406 438938 482448 439174
rect 482128 438854 482448 438938
rect 482128 438618 482170 438854
rect 482406 438618 482448 438854
rect 482128 438586 482448 438618
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 477008 399454 477328 399486
rect 477008 399218 477050 399454
rect 477286 399218 477328 399454
rect 477008 399134 477328 399218
rect 477008 398898 477050 399134
rect 477286 398898 477328 399134
rect 477008 398866 477328 398898
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 471888 346054 472208 346086
rect 471888 345818 471930 346054
rect 472166 345818 472208 346054
rect 471888 345734 472208 345818
rect 471888 345498 471930 345734
rect 472166 345498 472208 345734
rect 471888 345466 472208 345498
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 466768 306334 467088 306366
rect 466768 306098 466810 306334
rect 467046 306098 467088 306334
rect 466768 306014 467088 306098
rect 466768 305778 466810 306014
rect 467046 305778 467088 306014
rect 466768 305746 467088 305778
rect 461648 302614 461968 302646
rect 461648 302378 461690 302614
rect 461926 302378 461968 302614
rect 461648 302294 461968 302378
rect 461648 302058 461690 302294
rect 461926 302058 461968 302294
rect 461648 302026 461968 302058
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 456528 262894 456848 262926
rect 456528 262658 456570 262894
rect 456806 262658 456848 262894
rect 456528 262574 456848 262658
rect 456528 262338 456570 262574
rect 456806 262338 456848 262574
rect 456528 262306 456848 262338
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 451408 223174 451728 223206
rect 451408 222938 451450 223174
rect 451686 222938 451728 223174
rect 451408 222854 451728 222938
rect 451408 222618 451450 222854
rect 451686 222618 451728 222854
rect 451408 222586 451728 222618
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 446288 183454 446608 183486
rect 446288 183218 446330 183454
rect 446566 183218 446608 183454
rect 446288 183134 446608 183218
rect 446288 182898 446330 183134
rect 446566 182898 446608 183134
rect 446288 182866 446608 182898
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 441168 130054 441488 130086
rect 441168 129818 441210 130054
rect 441446 129818 441488 130054
rect 441168 129734 441488 129818
rect 441168 129498 441210 129734
rect 441446 129498 441488 129734
rect 441168 129466 441488 129498
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 436048 90334 436368 90366
rect 436048 90098 436090 90334
rect 436326 90098 436368 90334
rect 436048 90014 436368 90098
rect 436048 89778 436090 90014
rect 436326 89778 436368 90014
rect 436048 89746 436368 89778
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 430928 50614 431248 50646
rect 430928 50378 430970 50614
rect 431206 50378 431248 50614
rect 430928 50294 431248 50378
rect 430928 50058 430970 50294
rect 431206 50058 431248 50294
rect 430928 50026 431248 50058
rect 425808 46894 426128 46926
rect 425808 46658 425850 46894
rect 426086 46658 426128 46894
rect 425808 46574 426128 46658
rect 425808 46338 425850 46574
rect 426086 46338 426128 46574
rect 425808 46306 426128 46338
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 349008 22054 349328 22086
rect 349008 21818 349050 22054
rect 349286 21818 349328 22054
rect 349008 21734 349328 21818
rect 349008 21498 349050 21734
rect 349286 21498 349328 21734
rect 349008 21466 349328 21498
rect 379728 22054 380048 22086
rect 379728 21818 379770 22054
rect 380006 21818 380048 22054
rect 379728 21734 380048 21818
rect 379728 21498 379770 21734
rect 380006 21498 380048 21734
rect 379728 21466 380048 21498
rect 410448 22054 410768 22086
rect 410448 21818 410490 22054
rect 410726 21818 410768 22054
rect 410448 21734 410768 21818
rect 410448 21498 410490 21734
rect 410726 21498 410768 21734
rect 410448 21466 410768 21498
rect 343888 18334 344208 18366
rect 343888 18098 343930 18334
rect 344166 18098 344208 18334
rect 343888 18014 344208 18098
rect 343888 17778 343930 18014
rect 344166 17778 344208 18014
rect 343888 17746 344208 17778
rect 374608 18334 374928 18366
rect 374608 18098 374650 18334
rect 374886 18098 374928 18334
rect 374608 18014 374928 18098
rect 374608 17778 374650 18014
rect 374886 17778 374928 18014
rect 374608 17746 374928 17778
rect 405328 18334 405648 18366
rect 405328 18098 405370 18334
rect 405606 18098 405648 18334
rect 405328 18014 405648 18098
rect 405328 17778 405370 18014
rect 405606 17778 405648 18014
rect 405328 17746 405648 17778
rect 338768 14614 339088 14646
rect 338768 14378 338810 14614
rect 339046 14378 339088 14614
rect 338768 14294 339088 14378
rect 338768 14058 338810 14294
rect 339046 14058 339088 14294
rect 338768 14026 339088 14058
rect 369488 14614 369808 14646
rect 369488 14378 369530 14614
rect 369766 14378 369808 14614
rect 369488 14294 369808 14378
rect 369488 14058 369530 14294
rect 369766 14058 369808 14294
rect 369488 14026 369808 14058
rect 400208 14614 400528 14646
rect 400208 14378 400250 14614
rect 400486 14378 400528 14614
rect 400208 14294 400528 14378
rect 400208 14058 400250 14294
rect 400486 14058 400528 14294
rect 400208 14026 400528 14058
rect 333648 10894 333968 10926
rect 333648 10658 333690 10894
rect 333926 10658 333968 10894
rect 333648 10574 333968 10658
rect 333648 10338 333690 10574
rect 333926 10338 333968 10574
rect 333648 10306 333968 10338
rect 364368 10894 364688 10926
rect 364368 10658 364410 10894
rect 364646 10658 364688 10894
rect 364368 10574 364688 10658
rect 364368 10338 364410 10574
rect 364646 10338 364688 10574
rect 364368 10306 364688 10338
rect 395088 10894 395408 10926
rect 395088 10658 395130 10894
rect 395366 10658 395408 10894
rect 395088 10574 395408 10658
rect 395088 10338 395130 10574
rect 395366 10338 395408 10574
rect 395088 10306 395408 10338
rect 328528 7174 328848 7206
rect 328528 6938 328570 7174
rect 328806 6938 328848 7174
rect 328528 6854 328848 6938
rect 328528 6618 328570 6854
rect 328806 6618 328848 6854
rect 328528 6586 328848 6618
rect 359248 7174 359568 7206
rect 359248 6938 359290 7174
rect 359526 6938 359568 7174
rect 359248 6854 359568 6938
rect 359248 6618 359290 6854
rect 359526 6618 359568 6854
rect 359248 6586 359568 6618
rect 389968 7174 390288 7206
rect 389968 6938 390010 7174
rect 390246 6938 390288 7174
rect 389968 6854 390288 6938
rect 389968 6618 390010 6854
rect 390246 6618 390288 6854
rect 389968 6586 390288 6618
rect 420688 7174 421008 7206
rect 420688 6938 420730 7174
rect 420966 6938 421008 7174
rect 420688 6854 421008 6938
rect 420688 6618 420730 6854
rect 420966 6618 421008 6854
rect 420688 6586 421008 6618
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 -1306 330134 3479
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 -2266 333854 2988
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 -3226 337574 3479
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 -4186 341294 3479
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 -5146 345014 3479
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 -6106 348734 3479
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 -7066 352454 3479
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 3454 362414 3486
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 -1306 366134 3479
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 -2266 369854 2988
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 -3226 373574 3479
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 -4186 377294 3479
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 -5146 381014 3479
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 -6106 384734 2988
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 -7066 388454 3479
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 3454 398414 3486
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 -1306 402134 3479
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 -2266 405854 2988
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 -3226 409574 3479
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 -4186 413294 3479
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 -5146 417014 3479
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 -6106 420734 2988
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 -7066 424454 28938
rect 433794 39454 434414 74898
rect 437514 79174 438134 114618
rect 444954 122614 445574 158058
rect 448674 162334 449294 197778
rect 452394 202054 453014 237498
rect 459834 245494 460454 280938
rect 469794 291454 470414 326898
rect 473514 331174 474134 366618
rect 480954 374614 481574 410058
rect 484674 414334 485294 449778
rect 488394 454054 489014 489498
rect 495834 497494 496454 532938
rect 505794 543454 506414 578898
rect 507728 579454 508048 579486
rect 507728 579218 507770 579454
rect 508006 579218 508048 579454
rect 507728 579134 508048 579218
rect 507728 578898 507770 579134
rect 508006 578898 508048 579134
rect 507728 578866 508048 578898
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 502608 526054 502928 526086
rect 502608 525818 502650 526054
rect 502886 525818 502928 526054
rect 502608 525734 502928 525818
rect 502608 525498 502650 525734
rect 502886 525498 502928 525734
rect 502608 525466 502928 525498
rect 497488 522334 497808 522366
rect 497488 522098 497530 522334
rect 497766 522098 497808 522334
rect 497488 522014 497808 522098
rect 497488 521778 497530 522014
rect 497766 521778 497808 522014
rect 497488 521746 497808 521778
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 492368 482614 492688 482646
rect 492368 482378 492410 482614
rect 492646 482378 492688 482614
rect 492368 482294 492688 482378
rect 492368 482058 492410 482294
rect 492646 482058 492688 482294
rect 492368 482026 492688 482058
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 487248 442894 487568 442926
rect 487248 442658 487290 442894
rect 487526 442658 487568 442894
rect 487248 442574 487568 442658
rect 487248 442338 487290 442574
rect 487526 442338 487568 442574
rect 487248 442306 487568 442338
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 482128 403174 482448 403206
rect 482128 402938 482170 403174
rect 482406 402938 482448 403174
rect 482128 402854 482448 402938
rect 482128 402618 482170 402854
rect 482406 402618 482448 402854
rect 482128 402586 482448 402618
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 477008 363454 477328 363486
rect 477008 363218 477050 363454
rect 477286 363218 477328 363454
rect 477008 363134 477328 363218
rect 477008 362898 477050 363134
rect 477286 362898 477328 363134
rect 477008 362866 477328 362898
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 471888 310054 472208 310086
rect 471888 309818 471930 310054
rect 472166 309818 472208 310054
rect 471888 309734 472208 309818
rect 471888 309498 471930 309734
rect 472166 309498 472208 309734
rect 471888 309466 472208 309498
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 466768 270334 467088 270366
rect 466768 270098 466810 270334
rect 467046 270098 467088 270334
rect 466768 270014 467088 270098
rect 466768 269778 466810 270014
rect 467046 269778 467088 270014
rect 466768 269746 467088 269778
rect 461648 266614 461968 266646
rect 461648 266378 461690 266614
rect 461926 266378 461968 266614
rect 461648 266294 461968 266378
rect 461648 266058 461690 266294
rect 461926 266058 461968 266294
rect 461648 266026 461968 266058
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 456528 226894 456848 226926
rect 456528 226658 456570 226894
rect 456806 226658 456848 226894
rect 456528 226574 456848 226658
rect 456528 226338 456570 226574
rect 456806 226338 456848 226574
rect 456528 226306 456848 226338
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 451408 187174 451728 187206
rect 451408 186938 451450 187174
rect 451686 186938 451728 187174
rect 451408 186854 451728 186938
rect 451408 186618 451450 186854
rect 451686 186618 451728 186854
rect 451408 186586 451728 186618
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 446288 147454 446608 147486
rect 446288 147218 446330 147454
rect 446566 147218 446608 147454
rect 446288 147134 446608 147218
rect 446288 146898 446330 147134
rect 446566 146898 446608 147134
rect 446288 146866 446608 146898
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 441168 94054 441488 94086
rect 441168 93818 441210 94054
rect 441446 93818 441488 94054
rect 441168 93734 441488 93818
rect 441168 93498 441210 93734
rect 441446 93498 441488 93734
rect 441168 93466 441488 93498
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 436048 54334 436368 54366
rect 436048 54098 436090 54334
rect 436326 54098 436368 54334
rect 436048 54014 436368 54098
rect 436048 53778 436090 54014
rect 436326 53778 436368 54014
rect 436048 53746 436368 53778
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 430928 14614 431248 14646
rect 430928 14378 430970 14614
rect 431206 14378 431248 14614
rect 430928 14294 431248 14378
rect 430928 14058 430970 14294
rect 431206 14058 431248 14294
rect 430928 14026 431248 14058
rect 425808 10894 426128 10926
rect 425808 10658 425850 10894
rect 426086 10658 426128 10894
rect 425808 10574 426128 10658
rect 425808 10338 425850 10574
rect 426086 10338 426128 10574
rect 425808 10306 426128 10338
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 38898
rect 437514 43174 438134 78618
rect 444954 86614 445574 122058
rect 448674 126334 449294 161778
rect 452394 166054 453014 201498
rect 459834 209494 460454 244938
rect 469794 255454 470414 290898
rect 473514 295174 474134 330618
rect 480954 338614 481574 374058
rect 484674 378334 485294 413778
rect 488394 418054 489014 453498
rect 495834 461494 496454 496938
rect 505794 507454 506414 542898
rect 507728 543454 508048 543486
rect 507728 543218 507770 543454
rect 508006 543218 508048 543454
rect 507728 543134 508048 543218
rect 507728 542898 507770 543134
rect 508006 542898 508048 543134
rect 507728 542866 508048 542898
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 502608 490054 502928 490086
rect 502608 489818 502650 490054
rect 502886 489818 502928 490054
rect 502608 489734 502928 489818
rect 502608 489498 502650 489734
rect 502886 489498 502928 489734
rect 502608 489466 502928 489498
rect 497488 486334 497808 486366
rect 497488 486098 497530 486334
rect 497766 486098 497808 486334
rect 497488 486014 497808 486098
rect 497488 485778 497530 486014
rect 497766 485778 497808 486014
rect 497488 485746 497808 485778
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 492368 446614 492688 446646
rect 492368 446378 492410 446614
rect 492646 446378 492688 446614
rect 492368 446294 492688 446378
rect 492368 446058 492410 446294
rect 492646 446058 492688 446294
rect 492368 446026 492688 446058
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 487248 406894 487568 406926
rect 487248 406658 487290 406894
rect 487526 406658 487568 406894
rect 487248 406574 487568 406658
rect 487248 406338 487290 406574
rect 487526 406338 487568 406574
rect 487248 406306 487568 406338
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 482128 367174 482448 367206
rect 482128 366938 482170 367174
rect 482406 366938 482448 367174
rect 482128 366854 482448 366938
rect 482128 366618 482170 366854
rect 482406 366618 482448 366854
rect 482128 366586 482448 366618
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 477008 327454 477328 327486
rect 477008 327218 477050 327454
rect 477286 327218 477328 327454
rect 477008 327134 477328 327218
rect 477008 326898 477050 327134
rect 477286 326898 477328 327134
rect 477008 326866 477328 326898
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 471888 274054 472208 274086
rect 471888 273818 471930 274054
rect 472166 273818 472208 274054
rect 471888 273734 472208 273818
rect 471888 273498 471930 273734
rect 472166 273498 472208 273734
rect 471888 273466 472208 273498
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 466768 234334 467088 234366
rect 466768 234098 466810 234334
rect 467046 234098 467088 234334
rect 466768 234014 467088 234098
rect 466768 233778 466810 234014
rect 467046 233778 467088 234014
rect 466768 233746 467088 233778
rect 461648 230614 461968 230646
rect 461648 230378 461690 230614
rect 461926 230378 461968 230614
rect 461648 230294 461968 230378
rect 461648 230058 461690 230294
rect 461926 230058 461968 230294
rect 461648 230026 461968 230058
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 456528 190894 456848 190926
rect 456528 190658 456570 190894
rect 456806 190658 456848 190894
rect 456528 190574 456848 190658
rect 456528 190338 456570 190574
rect 456806 190338 456848 190574
rect 456528 190306 456848 190338
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 451408 151174 451728 151206
rect 451408 150938 451450 151174
rect 451686 150938 451728 151174
rect 451408 150854 451728 150938
rect 451408 150618 451450 150854
rect 451686 150618 451728 150854
rect 451408 150586 451728 150618
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 446288 111454 446608 111486
rect 446288 111218 446330 111454
rect 446566 111218 446608 111454
rect 446288 111134 446608 111218
rect 446288 110898 446330 111134
rect 446566 110898 446608 111134
rect 446288 110866 446608 110898
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 441168 58054 441488 58086
rect 441168 57818 441210 58054
rect 441446 57818 441488 58054
rect 441168 57734 441488 57818
rect 441168 57498 441210 57734
rect 441446 57498 441488 57734
rect 441168 57466 441488 57498
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 436048 18334 436368 18366
rect 436048 18098 436090 18334
rect 436326 18098 436368 18334
rect 436048 18014 436368 18098
rect 436048 17778 436090 18014
rect 436326 17778 436368 18014
rect 436048 17746 436368 17778
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 42618
rect 444954 50614 445574 86058
rect 448674 90334 449294 125778
rect 452394 130054 453014 165498
rect 459834 173494 460454 208938
rect 469794 219454 470414 254898
rect 473514 259174 474134 294618
rect 480954 302614 481574 338058
rect 484674 342334 485294 377778
rect 488394 382054 489014 417498
rect 495834 425494 496454 460938
rect 505794 471454 506414 506898
rect 507728 507454 508048 507486
rect 507728 507218 507770 507454
rect 508006 507218 508048 507454
rect 507728 507134 508048 507218
rect 507728 506898 507770 507134
rect 508006 506898 508048 507134
rect 507728 506866 508048 506898
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 502608 454054 502928 454086
rect 502608 453818 502650 454054
rect 502886 453818 502928 454054
rect 502608 453734 502928 453818
rect 502608 453498 502650 453734
rect 502886 453498 502928 453734
rect 502608 453466 502928 453498
rect 497488 450334 497808 450366
rect 497488 450098 497530 450334
rect 497766 450098 497808 450334
rect 497488 450014 497808 450098
rect 497488 449778 497530 450014
rect 497766 449778 497808 450014
rect 497488 449746 497808 449778
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 492368 410614 492688 410646
rect 492368 410378 492410 410614
rect 492646 410378 492688 410614
rect 492368 410294 492688 410378
rect 492368 410058 492410 410294
rect 492646 410058 492688 410294
rect 492368 410026 492688 410058
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 487248 370894 487568 370926
rect 487248 370658 487290 370894
rect 487526 370658 487568 370894
rect 487248 370574 487568 370658
rect 487248 370338 487290 370574
rect 487526 370338 487568 370574
rect 487248 370306 487568 370338
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 482128 331174 482448 331206
rect 482128 330938 482170 331174
rect 482406 330938 482448 331174
rect 482128 330854 482448 330938
rect 482128 330618 482170 330854
rect 482406 330618 482448 330854
rect 482128 330586 482448 330618
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 477008 291454 477328 291486
rect 477008 291218 477050 291454
rect 477286 291218 477328 291454
rect 477008 291134 477328 291218
rect 477008 290898 477050 291134
rect 477286 290898 477328 291134
rect 477008 290866 477328 290898
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 471888 238054 472208 238086
rect 471888 237818 471930 238054
rect 472166 237818 472208 238054
rect 471888 237734 472208 237818
rect 471888 237498 471930 237734
rect 472166 237498 472208 237734
rect 471888 237466 472208 237498
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 466768 198334 467088 198366
rect 466768 198098 466810 198334
rect 467046 198098 467088 198334
rect 466768 198014 467088 198098
rect 466768 197778 466810 198014
rect 467046 197778 467088 198014
rect 466768 197746 467088 197778
rect 461648 194614 461968 194646
rect 461648 194378 461690 194614
rect 461926 194378 461968 194614
rect 461648 194294 461968 194378
rect 461648 194058 461690 194294
rect 461926 194058 461968 194294
rect 461648 194026 461968 194058
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 456528 154894 456848 154926
rect 456528 154658 456570 154894
rect 456806 154658 456848 154894
rect 456528 154574 456848 154658
rect 456528 154338 456570 154574
rect 456806 154338 456848 154574
rect 456528 154306 456848 154338
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 451408 115174 451728 115206
rect 451408 114938 451450 115174
rect 451686 114938 451728 115174
rect 451408 114854 451728 114938
rect 451408 114618 451450 114854
rect 451686 114618 451728 114854
rect 451408 114586 451728 114618
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 446288 75454 446608 75486
rect 446288 75218 446330 75454
rect 446566 75218 446608 75454
rect 446288 75134 446608 75218
rect 446288 74898 446330 75134
rect 446566 74898 446608 75134
rect 446288 74866 446608 74898
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 441168 22054 441488 22086
rect 441168 21818 441210 22054
rect 441446 21818 441488 22054
rect 441168 21734 441488 21818
rect 441168 21498 441210 21734
rect 441446 21498 441488 21734
rect 441168 21466 441488 21498
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 444954 14614 445574 50058
rect 448674 54334 449294 89778
rect 452394 94054 453014 129498
rect 459834 137494 460454 172938
rect 469794 183454 470414 218898
rect 473514 223174 474134 258618
rect 480954 266614 481574 302058
rect 484674 306334 485294 341778
rect 488394 346054 489014 381498
rect 495834 389494 496454 424938
rect 505794 435454 506414 470898
rect 507728 471454 508048 471486
rect 507728 471218 507770 471454
rect 508006 471218 508048 471454
rect 507728 471134 508048 471218
rect 507728 470898 507770 471134
rect 508006 470898 508048 471134
rect 507728 470866 508048 470898
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 502608 418054 502928 418086
rect 502608 417818 502650 418054
rect 502886 417818 502928 418054
rect 502608 417734 502928 417818
rect 502608 417498 502650 417734
rect 502886 417498 502928 417734
rect 502608 417466 502928 417498
rect 497488 414334 497808 414366
rect 497488 414098 497530 414334
rect 497766 414098 497808 414334
rect 497488 414014 497808 414098
rect 497488 413778 497530 414014
rect 497766 413778 497808 414014
rect 497488 413746 497808 413778
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 492368 374614 492688 374646
rect 492368 374378 492410 374614
rect 492646 374378 492688 374614
rect 492368 374294 492688 374378
rect 492368 374058 492410 374294
rect 492646 374058 492688 374294
rect 492368 374026 492688 374058
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 487248 334894 487568 334926
rect 487248 334658 487290 334894
rect 487526 334658 487568 334894
rect 487248 334574 487568 334658
rect 487248 334338 487290 334574
rect 487526 334338 487568 334574
rect 487248 334306 487568 334338
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 482128 295174 482448 295206
rect 482128 294938 482170 295174
rect 482406 294938 482448 295174
rect 482128 294854 482448 294938
rect 482128 294618 482170 294854
rect 482406 294618 482448 294854
rect 482128 294586 482448 294618
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 477008 255454 477328 255486
rect 477008 255218 477050 255454
rect 477286 255218 477328 255454
rect 477008 255134 477328 255218
rect 477008 254898 477050 255134
rect 477286 254898 477328 255134
rect 477008 254866 477328 254898
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 471888 202054 472208 202086
rect 471888 201818 471930 202054
rect 472166 201818 472208 202054
rect 471888 201734 472208 201818
rect 471888 201498 471930 201734
rect 472166 201498 472208 201734
rect 471888 201466 472208 201498
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 466768 162334 467088 162366
rect 466768 162098 466810 162334
rect 467046 162098 467088 162334
rect 466768 162014 467088 162098
rect 466768 161778 466810 162014
rect 467046 161778 467088 162014
rect 466768 161746 467088 161778
rect 461648 158614 461968 158646
rect 461648 158378 461690 158614
rect 461926 158378 461968 158614
rect 461648 158294 461968 158378
rect 461648 158058 461690 158294
rect 461926 158058 461968 158294
rect 461648 158026 461968 158058
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 456528 118894 456848 118926
rect 456528 118658 456570 118894
rect 456806 118658 456848 118894
rect 456528 118574 456848 118658
rect 456528 118338 456570 118574
rect 456806 118338 456848 118574
rect 456528 118306 456848 118338
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 451408 79174 451728 79206
rect 451408 78938 451450 79174
rect 451686 78938 451728 79174
rect 451408 78854 451728 78938
rect 451408 78618 451450 78854
rect 451686 78618 451728 78854
rect 451408 78586 451728 78618
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 446288 39454 446608 39486
rect 446288 39218 446330 39454
rect 446566 39218 446608 39454
rect 446288 39134 446608 39218
rect 446288 38898 446330 39134
rect 446566 38898 446608 39134
rect 446288 38866 446608 38898
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 -2266 441854 2988
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 53778
rect 452394 58054 453014 93498
rect 459834 101494 460454 136938
rect 469794 147454 470414 182898
rect 473514 187174 474134 222618
rect 480954 230614 481574 266058
rect 484674 270334 485294 305778
rect 488394 310054 489014 345498
rect 495834 353494 496454 388938
rect 505794 399454 506414 434898
rect 507728 435454 508048 435486
rect 507728 435218 507770 435454
rect 508006 435218 508048 435454
rect 507728 435134 508048 435218
rect 507728 434898 507770 435134
rect 508006 434898 508048 435134
rect 507728 434866 508048 434898
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 502608 382054 502928 382086
rect 502608 381818 502650 382054
rect 502886 381818 502928 382054
rect 502608 381734 502928 381818
rect 502608 381498 502650 381734
rect 502886 381498 502928 381734
rect 502608 381466 502928 381498
rect 497488 378334 497808 378366
rect 497488 378098 497530 378334
rect 497766 378098 497808 378334
rect 497488 378014 497808 378098
rect 497488 377778 497530 378014
rect 497766 377778 497808 378014
rect 497488 377746 497808 377778
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 492368 338614 492688 338646
rect 492368 338378 492410 338614
rect 492646 338378 492688 338614
rect 492368 338294 492688 338378
rect 492368 338058 492410 338294
rect 492646 338058 492688 338294
rect 492368 338026 492688 338058
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 487248 298894 487568 298926
rect 487248 298658 487290 298894
rect 487526 298658 487568 298894
rect 487248 298574 487568 298658
rect 487248 298338 487290 298574
rect 487526 298338 487568 298574
rect 487248 298306 487568 298338
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 482128 259174 482448 259206
rect 482128 258938 482170 259174
rect 482406 258938 482448 259174
rect 482128 258854 482448 258938
rect 482128 258618 482170 258854
rect 482406 258618 482448 258854
rect 482128 258586 482448 258618
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 477008 219454 477328 219486
rect 477008 219218 477050 219454
rect 477286 219218 477328 219454
rect 477008 219134 477328 219218
rect 477008 218898 477050 219134
rect 477286 218898 477328 219134
rect 477008 218866 477328 218898
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 471888 166054 472208 166086
rect 471888 165818 471930 166054
rect 472166 165818 472208 166054
rect 471888 165734 472208 165818
rect 471888 165498 471930 165734
rect 472166 165498 472208 165734
rect 471888 165466 472208 165498
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 466768 126334 467088 126366
rect 466768 126098 466810 126334
rect 467046 126098 467088 126334
rect 466768 126014 467088 126098
rect 466768 125778 466810 126014
rect 467046 125778 467088 126014
rect 466768 125746 467088 125778
rect 461648 122614 461968 122646
rect 461648 122378 461690 122614
rect 461926 122378 461968 122614
rect 461648 122294 461968 122378
rect 461648 122058 461690 122294
rect 461926 122058 461968 122294
rect 461648 122026 461968 122058
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 456528 82894 456848 82926
rect 456528 82658 456570 82894
rect 456806 82658 456848 82894
rect 456528 82574 456848 82658
rect 456528 82338 456570 82574
rect 456806 82338 456848 82574
rect 456528 82306 456848 82338
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 451408 43174 451728 43206
rect 451408 42938 451450 43174
rect 451686 42938 451728 43174
rect 451408 42854 451728 42938
rect 451408 42618 451450 42854
rect 451686 42618 451728 42854
rect 451408 42586 451728 42618
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 452394 22054 453014 57498
rect 459834 65494 460454 100938
rect 469794 111454 470414 146898
rect 473514 151174 474134 186618
rect 480954 194614 481574 230058
rect 484674 234334 485294 269778
rect 488394 274054 489014 309498
rect 495834 317494 496454 352938
rect 505794 363454 506414 398898
rect 507728 399454 508048 399486
rect 507728 399218 507770 399454
rect 508006 399218 508048 399454
rect 507728 399134 508048 399218
rect 507728 398898 507770 399134
rect 508006 398898 508048 399134
rect 507728 398866 508048 398898
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 502608 346054 502928 346086
rect 502608 345818 502650 346054
rect 502886 345818 502928 346054
rect 502608 345734 502928 345818
rect 502608 345498 502650 345734
rect 502886 345498 502928 345734
rect 502608 345466 502928 345498
rect 497488 342334 497808 342366
rect 497488 342098 497530 342334
rect 497766 342098 497808 342334
rect 497488 342014 497808 342098
rect 497488 341778 497530 342014
rect 497766 341778 497808 342014
rect 497488 341746 497808 341778
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 492368 302614 492688 302646
rect 492368 302378 492410 302614
rect 492646 302378 492688 302614
rect 492368 302294 492688 302378
rect 492368 302058 492410 302294
rect 492646 302058 492688 302294
rect 492368 302026 492688 302058
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 487248 262894 487568 262926
rect 487248 262658 487290 262894
rect 487526 262658 487568 262894
rect 487248 262574 487568 262658
rect 487248 262338 487290 262574
rect 487526 262338 487568 262574
rect 487248 262306 487568 262338
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 482128 223174 482448 223206
rect 482128 222938 482170 223174
rect 482406 222938 482448 223174
rect 482128 222854 482448 222938
rect 482128 222618 482170 222854
rect 482406 222618 482448 222854
rect 482128 222586 482448 222618
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 477008 183454 477328 183486
rect 477008 183218 477050 183454
rect 477286 183218 477328 183454
rect 477008 183134 477328 183218
rect 477008 182898 477050 183134
rect 477286 182898 477328 183134
rect 477008 182866 477328 182898
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 471888 130054 472208 130086
rect 471888 129818 471930 130054
rect 472166 129818 472208 130054
rect 471888 129734 472208 129818
rect 471888 129498 471930 129734
rect 472166 129498 472208 129734
rect 471888 129466 472208 129498
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 466768 90334 467088 90366
rect 466768 90098 466810 90334
rect 467046 90098 467088 90334
rect 466768 90014 467088 90098
rect 466768 89778 466810 90014
rect 467046 89778 467088 90014
rect 466768 89746 467088 89778
rect 461648 86614 461968 86646
rect 461648 86378 461690 86614
rect 461926 86378 461968 86614
rect 461648 86294 461968 86378
rect 461648 86058 461690 86294
rect 461926 86058 461968 86294
rect 461648 86026 461968 86058
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 456528 46894 456848 46926
rect 456528 46658 456570 46894
rect 456806 46658 456848 46894
rect 456528 46574 456848 46658
rect 456528 46338 456570 46574
rect 456806 46338 456848 46574
rect 456528 46306 456848 46338
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 451408 7174 451728 7206
rect 451408 6938 451450 7174
rect 451686 6938 451728 7174
rect 451408 6854 451728 6938
rect 451408 6618 451450 6854
rect 451686 6618 451728 6854
rect 451408 6586 451728 6618
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 -5146 453014 21498
rect 459834 29494 460454 64938
rect 469794 75454 470414 110898
rect 473514 115174 474134 150618
rect 480954 158614 481574 194058
rect 484674 198334 485294 233778
rect 488394 238054 489014 273498
rect 495834 281494 496454 316938
rect 505794 327454 506414 362898
rect 507728 363454 508048 363486
rect 507728 363218 507770 363454
rect 508006 363218 508048 363454
rect 507728 363134 508048 363218
rect 507728 362898 507770 363134
rect 508006 362898 508048 363134
rect 507728 362866 508048 362898
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 502608 310054 502928 310086
rect 502608 309818 502650 310054
rect 502886 309818 502928 310054
rect 502608 309734 502928 309818
rect 502608 309498 502650 309734
rect 502886 309498 502928 309734
rect 502608 309466 502928 309498
rect 497488 306334 497808 306366
rect 497488 306098 497530 306334
rect 497766 306098 497808 306334
rect 497488 306014 497808 306098
rect 497488 305778 497530 306014
rect 497766 305778 497808 306014
rect 497488 305746 497808 305778
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 492368 266614 492688 266646
rect 492368 266378 492410 266614
rect 492646 266378 492688 266614
rect 492368 266294 492688 266378
rect 492368 266058 492410 266294
rect 492646 266058 492688 266294
rect 492368 266026 492688 266058
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 487248 226894 487568 226926
rect 487248 226658 487290 226894
rect 487526 226658 487568 226894
rect 487248 226574 487568 226658
rect 487248 226338 487290 226574
rect 487526 226338 487568 226574
rect 487248 226306 487568 226338
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 482128 187174 482448 187206
rect 482128 186938 482170 187174
rect 482406 186938 482448 187174
rect 482128 186854 482448 186938
rect 482128 186618 482170 186854
rect 482406 186618 482448 186854
rect 482128 186586 482448 186618
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 477008 147454 477328 147486
rect 477008 147218 477050 147454
rect 477286 147218 477328 147454
rect 477008 147134 477328 147218
rect 477008 146898 477050 147134
rect 477286 146898 477328 147134
rect 477008 146866 477328 146898
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 471888 94054 472208 94086
rect 471888 93818 471930 94054
rect 472166 93818 472208 94054
rect 471888 93734 472208 93818
rect 471888 93498 471930 93734
rect 472166 93498 472208 93734
rect 471888 93466 472208 93498
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 466768 54334 467088 54366
rect 466768 54098 466810 54334
rect 467046 54098 467088 54334
rect 466768 54014 467088 54098
rect 466768 53778 466810 54014
rect 467046 53778 467088 54014
rect 466768 53746 467088 53778
rect 461648 50614 461968 50646
rect 461648 50378 461690 50614
rect 461926 50378 461968 50614
rect 461648 50294 461968 50378
rect 461648 50058 461690 50294
rect 461926 50058 461968 50294
rect 461648 50026 461968 50058
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 456528 10894 456848 10926
rect 456528 10658 456570 10894
rect 456806 10658 456848 10894
rect 456528 10574 456848 10658
rect 456528 10338 456570 10574
rect 456806 10338 456848 10574
rect 456528 10306 456848 10338
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 -6106 456734 2988
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 -7066 460454 28938
rect 469794 39454 470414 74898
rect 473514 79174 474134 114618
rect 480954 122614 481574 158058
rect 484674 162334 485294 197778
rect 488394 202054 489014 237498
rect 495834 245494 496454 280938
rect 505794 291454 506414 326898
rect 507728 327454 508048 327486
rect 507728 327218 507770 327454
rect 508006 327218 508048 327454
rect 507728 327134 508048 327218
rect 507728 326898 507770 327134
rect 508006 326898 508048 327134
rect 507728 326866 508048 326898
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 502608 274054 502928 274086
rect 502608 273818 502650 274054
rect 502886 273818 502928 274054
rect 502608 273734 502928 273818
rect 502608 273498 502650 273734
rect 502886 273498 502928 273734
rect 502608 273466 502928 273498
rect 497488 270334 497808 270366
rect 497488 270098 497530 270334
rect 497766 270098 497808 270334
rect 497488 270014 497808 270098
rect 497488 269778 497530 270014
rect 497766 269778 497808 270014
rect 497488 269746 497808 269778
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 492368 230614 492688 230646
rect 492368 230378 492410 230614
rect 492646 230378 492688 230614
rect 492368 230294 492688 230378
rect 492368 230058 492410 230294
rect 492646 230058 492688 230294
rect 492368 230026 492688 230058
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 487248 190894 487568 190926
rect 487248 190658 487290 190894
rect 487526 190658 487568 190894
rect 487248 190574 487568 190658
rect 487248 190338 487290 190574
rect 487526 190338 487568 190574
rect 487248 190306 487568 190338
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 482128 151174 482448 151206
rect 482128 150938 482170 151174
rect 482406 150938 482448 151174
rect 482128 150854 482448 150938
rect 482128 150618 482170 150854
rect 482406 150618 482448 150854
rect 482128 150586 482448 150618
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 477008 111454 477328 111486
rect 477008 111218 477050 111454
rect 477286 111218 477328 111454
rect 477008 111134 477328 111218
rect 477008 110898 477050 111134
rect 477286 110898 477328 111134
rect 477008 110866 477328 110898
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 471888 58054 472208 58086
rect 471888 57818 471930 58054
rect 472166 57818 472208 58054
rect 471888 57734 472208 57818
rect 471888 57498 471930 57734
rect 472166 57498 472208 57734
rect 471888 57466 472208 57498
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 466768 18334 467088 18366
rect 466768 18098 466810 18334
rect 467046 18098 467088 18334
rect 466768 18014 467088 18098
rect 466768 17778 466810 18014
rect 467046 17778 467088 18014
rect 466768 17746 467088 17778
rect 461648 14614 461968 14646
rect 461648 14378 461690 14614
rect 461926 14378 461968 14614
rect 461648 14294 461968 14378
rect 461648 14058 461690 14294
rect 461926 14058 461968 14294
rect 461648 14026 461968 14058
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 3454 470414 38898
rect 473514 43174 474134 78618
rect 480954 86614 481574 122058
rect 484674 126334 485294 161778
rect 488394 166054 489014 201498
rect 495834 209494 496454 244938
rect 505794 255454 506414 290898
rect 507728 291454 508048 291486
rect 507728 291218 507770 291454
rect 508006 291218 508048 291454
rect 507728 291134 508048 291218
rect 507728 290898 507770 291134
rect 508006 290898 508048 291134
rect 507728 290866 508048 290898
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 502608 238054 502928 238086
rect 502608 237818 502650 238054
rect 502886 237818 502928 238054
rect 502608 237734 502928 237818
rect 502608 237498 502650 237734
rect 502886 237498 502928 237734
rect 502608 237466 502928 237498
rect 497488 234334 497808 234366
rect 497488 234098 497530 234334
rect 497766 234098 497808 234334
rect 497488 234014 497808 234098
rect 497488 233778 497530 234014
rect 497766 233778 497808 234014
rect 497488 233746 497808 233778
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 492368 194614 492688 194646
rect 492368 194378 492410 194614
rect 492646 194378 492688 194614
rect 492368 194294 492688 194378
rect 492368 194058 492410 194294
rect 492646 194058 492688 194294
rect 492368 194026 492688 194058
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 487248 154894 487568 154926
rect 487248 154658 487290 154894
rect 487526 154658 487568 154894
rect 487248 154574 487568 154658
rect 487248 154338 487290 154574
rect 487526 154338 487568 154574
rect 487248 154306 487568 154338
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 482128 115174 482448 115206
rect 482128 114938 482170 115174
rect 482406 114938 482448 115174
rect 482128 114854 482448 114938
rect 482128 114618 482170 114854
rect 482406 114618 482448 114854
rect 482128 114586 482448 114618
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 477008 75454 477328 75486
rect 477008 75218 477050 75454
rect 477286 75218 477328 75454
rect 477008 75134 477328 75218
rect 477008 74898 477050 75134
rect 477286 74898 477328 75134
rect 477008 74866 477328 74898
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 471888 22054 472208 22086
rect 471888 21818 471930 22054
rect 472166 21818 472208 22054
rect 471888 21734 472208 21818
rect 471888 21498 471930 21734
rect 472166 21498 472208 21734
rect 471888 21466 472208 21498
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 42618
rect 480954 50614 481574 86058
rect 484674 90334 485294 125778
rect 488394 130054 489014 165498
rect 495834 173494 496454 208938
rect 505794 219454 506414 254898
rect 507728 255454 508048 255486
rect 507728 255218 507770 255454
rect 508006 255218 508048 255454
rect 507728 255134 508048 255218
rect 507728 254898 507770 255134
rect 508006 254898 508048 255134
rect 507728 254866 508048 254898
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 502608 202054 502928 202086
rect 502608 201818 502650 202054
rect 502886 201818 502928 202054
rect 502608 201734 502928 201818
rect 502608 201498 502650 201734
rect 502886 201498 502928 201734
rect 502608 201466 502928 201498
rect 497488 198334 497808 198366
rect 497488 198098 497530 198334
rect 497766 198098 497808 198334
rect 497488 198014 497808 198098
rect 497488 197778 497530 198014
rect 497766 197778 497808 198014
rect 497488 197746 497808 197778
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 492368 158614 492688 158646
rect 492368 158378 492410 158614
rect 492646 158378 492688 158614
rect 492368 158294 492688 158378
rect 492368 158058 492410 158294
rect 492646 158058 492688 158294
rect 492368 158026 492688 158058
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 487248 118894 487568 118926
rect 487248 118658 487290 118894
rect 487526 118658 487568 118894
rect 487248 118574 487568 118658
rect 487248 118338 487290 118574
rect 487526 118338 487568 118574
rect 487248 118306 487568 118338
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 482128 79174 482448 79206
rect 482128 78938 482170 79174
rect 482406 78938 482448 79174
rect 482128 78854 482448 78938
rect 482128 78618 482170 78854
rect 482406 78618 482448 78854
rect 482128 78586 482448 78618
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 477008 39454 477328 39486
rect 477008 39218 477050 39454
rect 477286 39218 477328 39454
rect 477008 39134 477328 39218
rect 477008 38898 477050 39134
rect 477286 38898 477328 39134
rect 477008 38866 477328 38898
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 480954 14614 481574 50058
rect 484674 54334 485294 89778
rect 488394 94054 489014 129498
rect 495834 137494 496454 172938
rect 505794 183454 506414 218898
rect 507728 219454 508048 219486
rect 507728 219218 507770 219454
rect 508006 219218 508048 219454
rect 507728 219134 508048 219218
rect 507728 218898 507770 219134
rect 508006 218898 508048 219134
rect 507728 218866 508048 218898
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 502608 166054 502928 166086
rect 502608 165818 502650 166054
rect 502886 165818 502928 166054
rect 502608 165734 502928 165818
rect 502608 165498 502650 165734
rect 502886 165498 502928 165734
rect 502608 165466 502928 165498
rect 497488 162334 497808 162366
rect 497488 162098 497530 162334
rect 497766 162098 497808 162334
rect 497488 162014 497808 162098
rect 497488 161778 497530 162014
rect 497766 161778 497808 162014
rect 497488 161746 497808 161778
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 492368 122614 492688 122646
rect 492368 122378 492410 122614
rect 492646 122378 492688 122614
rect 492368 122294 492688 122378
rect 492368 122058 492410 122294
rect 492646 122058 492688 122294
rect 492368 122026 492688 122058
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 487248 82894 487568 82926
rect 487248 82658 487290 82894
rect 487526 82658 487568 82894
rect 487248 82574 487568 82658
rect 487248 82338 487290 82574
rect 487526 82338 487568 82574
rect 487248 82306 487568 82338
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 482128 43174 482448 43206
rect 482128 42938 482170 43174
rect 482406 42938 482448 43174
rect 482128 42854 482448 42938
rect 482128 42618 482170 42854
rect 482406 42618 482448 42854
rect 482128 42586 482448 42618
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 -2266 477854 2988
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 -3226 481574 14058
rect 484674 18334 485294 53778
rect 488394 58054 489014 93498
rect 495834 101494 496454 136938
rect 505794 147454 506414 182898
rect 507728 183454 508048 183486
rect 507728 183218 507770 183454
rect 508006 183218 508048 183454
rect 507728 183134 508048 183218
rect 507728 182898 507770 183134
rect 508006 182898 508048 183134
rect 507728 182866 508048 182898
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 502608 130054 502928 130086
rect 502608 129818 502650 130054
rect 502886 129818 502928 130054
rect 502608 129734 502928 129818
rect 502608 129498 502650 129734
rect 502886 129498 502928 129734
rect 502608 129466 502928 129498
rect 497488 126334 497808 126366
rect 497488 126098 497530 126334
rect 497766 126098 497808 126334
rect 497488 126014 497808 126098
rect 497488 125778 497530 126014
rect 497766 125778 497808 126014
rect 497488 125746 497808 125778
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 492368 86614 492688 86646
rect 492368 86378 492410 86614
rect 492646 86378 492688 86614
rect 492368 86294 492688 86378
rect 492368 86058 492410 86294
rect 492646 86058 492688 86294
rect 492368 86026 492688 86058
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 487248 46894 487568 46926
rect 487248 46658 487290 46894
rect 487526 46658 487568 46894
rect 487248 46574 487568 46658
rect 487248 46338 487290 46574
rect 487526 46338 487568 46574
rect 487248 46306 487568 46338
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 482128 7174 482448 7206
rect 482128 6938 482170 7174
rect 482406 6938 482448 7174
rect 482128 6854 482448 6938
rect 482128 6618 482170 6854
rect 482406 6618 482448 6854
rect 482128 6586 482448 6618
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 -4186 485294 17778
rect 488394 22054 489014 57498
rect 495834 65494 496454 100938
rect 505794 111454 506414 146898
rect 507728 147454 508048 147486
rect 507728 147218 507770 147454
rect 508006 147218 508048 147454
rect 507728 147134 508048 147218
rect 507728 146898 507770 147134
rect 508006 146898 508048 147134
rect 507728 146866 508048 146898
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 502608 94054 502928 94086
rect 502608 93818 502650 94054
rect 502886 93818 502928 94054
rect 502608 93734 502928 93818
rect 502608 93498 502650 93734
rect 502886 93498 502928 93734
rect 502608 93466 502928 93498
rect 497488 90334 497808 90366
rect 497488 90098 497530 90334
rect 497766 90098 497808 90334
rect 497488 90014 497808 90098
rect 497488 89778 497530 90014
rect 497766 89778 497808 90014
rect 497488 89746 497808 89778
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 492368 50614 492688 50646
rect 492368 50378 492410 50614
rect 492646 50378 492688 50614
rect 492368 50294 492688 50378
rect 492368 50058 492410 50294
rect 492646 50058 492688 50294
rect 492368 50026 492688 50058
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 487248 10894 487568 10926
rect 487248 10658 487290 10894
rect 487526 10658 487568 10894
rect 487248 10574 487568 10658
rect 487248 10338 487290 10574
rect 487526 10338 487568 10574
rect 487248 10306 487568 10338
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 -5146 489014 21498
rect 495834 29494 496454 64938
rect 505794 75454 506414 110898
rect 507728 111454 508048 111486
rect 507728 111218 507770 111454
rect 508006 111218 508048 111454
rect 507728 111134 508048 111218
rect 507728 110898 507770 111134
rect 508006 110898 508048 111134
rect 507728 110866 508048 110898
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 502608 58054 502928 58086
rect 502608 57818 502650 58054
rect 502886 57818 502928 58054
rect 502608 57734 502928 57818
rect 502608 57498 502650 57734
rect 502886 57498 502928 57734
rect 502608 57466 502928 57498
rect 497488 54334 497808 54366
rect 497488 54098 497530 54334
rect 497766 54098 497808 54334
rect 497488 54014 497808 54098
rect 497488 53778 497530 54014
rect 497766 53778 497808 54014
rect 497488 53746 497808 53778
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 492368 14614 492688 14646
rect 492368 14378 492410 14614
rect 492646 14378 492688 14614
rect 492368 14294 492688 14378
rect 492368 14058 492410 14294
rect 492646 14058 492688 14294
rect 492368 14026 492688 14058
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 -6106 492734 2988
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 -7066 496454 28938
rect 505794 39454 506414 74898
rect 507728 75454 508048 75486
rect 507728 75218 507770 75454
rect 508006 75218 508048 75454
rect 507728 75134 508048 75218
rect 507728 74898 507770 75134
rect 508006 74898 508048 75134
rect 507728 74866 508048 74898
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 502608 22054 502928 22086
rect 502608 21818 502650 22054
rect 502886 21818 502928 22054
rect 502608 21734 502928 21818
rect 502608 21498 502650 21734
rect 502886 21498 502928 21734
rect 502608 21466 502928 21498
rect 497488 18334 497808 18366
rect 497488 18098 497530 18334
rect 497766 18098 497808 18334
rect 497488 18014 497808 18098
rect 497488 17778 497530 18014
rect 497766 17778 497808 18014
rect 497488 17746 497808 17778
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 3454 506414 38898
rect 507728 39454 508048 39486
rect 507728 39218 507770 39454
rect 508006 39218 508048 39454
rect 507728 39134 508048 39218
rect 507728 38898 507770 39134
rect 508006 38898 508048 39134
rect 507728 38866 508048 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 514155 644060 514221 644061
rect 514155 643996 514156 644060
rect 514220 643996 514221 644060
rect 514155 643995 514221 643996
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 514158 587077 514218 643995
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 514155 587076 514221 587077
rect 514155 587012 514156 587076
rect 514220 587012 514221 587076
rect 514155 587011 514221 587012
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 514155 537844 514221 537845
rect 514155 537780 514156 537844
rect 514220 537780 514221 537844
rect 514155 537779 514221 537780
rect 514158 527237 514218 537779
rect 514155 527236 514221 527237
rect 514155 527172 514156 527236
rect 514220 527172 514221 527236
rect 514155 527171 514221 527172
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 514155 497316 514221 497317
rect 514155 497252 514156 497316
rect 514220 497252 514221 497316
rect 514155 497251 514221 497252
rect 514158 484669 514218 497251
rect 514155 484668 514221 484669
rect 514155 484604 514156 484668
rect 514220 484604 514221 484668
rect 514155 484603 514221 484604
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 514339 467396 514405 467397
rect 514339 467332 514340 467396
rect 514404 467332 514405 467396
rect 514339 467331 514405 467332
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 514155 437476 514221 437477
rect 514155 437412 514156 437476
rect 514220 437412 514221 437476
rect 514155 437411 514221 437412
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 514158 378453 514218 437411
rect 514342 431629 514402 467331
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 514339 431628 514405 431629
rect 514339 431564 514340 431628
rect 514404 431564 514405 431628
rect 514339 431563 514405 431564
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 514339 407556 514405 407557
rect 514339 407492 514340 407556
rect 514404 407492 514405 407556
rect 514339 407491 514405 407492
rect 514155 378452 514221 378453
rect 514155 378388 514156 378452
rect 514220 378388 514221 378452
rect 514155 378387 514221 378388
rect 514155 377636 514221 377637
rect 514155 377572 514156 377636
rect 514220 377572 514221 377636
rect 514155 377571 514221 377572
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 514158 272237 514218 377571
rect 514342 325277 514402 407491
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 514339 325276 514405 325277
rect 514339 325212 514340 325276
rect 514404 325212 514405 325276
rect 514339 325211 514405 325212
rect 514339 317796 514405 317797
rect 514339 317732 514340 317796
rect 514404 317732 514405 317796
rect 514339 317731 514405 317732
rect 514155 272236 514221 272237
rect 514155 272172 514156 272236
rect 514220 272172 514221 272236
rect 514155 272171 514221 272172
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 514155 257956 514221 257957
rect 514155 257892 514156 257956
rect 514220 257892 514221 257956
rect 514155 257891 514221 257892
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 514158 112845 514218 257891
rect 514342 192541 514402 317731
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 514339 192540 514405 192541
rect 514339 192476 514340 192540
rect 514404 192476 514405 192540
rect 514339 192475 514405 192476
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 514155 112844 514221 112845
rect 514155 112780 514156 112844
rect 514220 112780 514221 112844
rect 514155 112779 514221 112780
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 580211 602308 580277 602309
rect 580211 602244 580212 602308
rect 580276 602244 580277 602308
rect 580211 602243 580277 602244
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 580214 205733 580274 602243
rect 580395 591020 580461 591021
rect 580395 590956 580396 591020
rect 580460 590956 580461 591020
rect 580395 590955 580461 590956
rect 580398 557157 580458 590955
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 580395 557156 580461 557157
rect 580395 557092 580396 557156
rect 580460 557092 580461 557156
rect 580395 557091 580461 557092
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 580395 219060 580461 219061
rect 580395 218996 580396 219060
rect 580460 218996 580461 219060
rect 580395 218995 580461 218996
rect 580211 205732 580277 205733
rect 580211 205668 580212 205732
rect 580276 205668 580277 205732
rect 580211 205667 580277 205668
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 580211 179212 580277 179213
rect 580211 179148 580212 179212
rect 580276 179148 580277 179212
rect 580211 179147 580277 179148
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 580214 138277 580274 179147
rect 580398 168197 580458 218995
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 580395 168196 580461 168197
rect 580395 168132 580396 168196
rect 580460 168132 580461 168196
rect 580395 168131 580461 168132
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 580395 139364 580461 139365
rect 580395 139300 580396 139364
rect 580460 139300 580461 139364
rect 580395 139299 580461 139300
rect 580211 138276 580277 138277
rect 580211 138212 580212 138276
rect 580276 138212 580277 138276
rect 580211 138211 580277 138212
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 580398 108357 580458 139299
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 580395 108356 580461 108357
rect 580395 108292 580396 108356
rect 580460 108292 580461 108356
rect 580395 108291 580461 108292
rect 580211 99516 580277 99517
rect 580211 99452 580212 99516
rect 580276 99452 580277 99516
rect 580211 99451 580277 99452
rect 580214 78437 580274 99451
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 580211 78436 580277 78437
rect 580211 78372 580212 78436
rect 580276 78372 580277 78436
rect 580211 78371 580277 78372
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 580211 59668 580277 59669
rect 580211 59604 580212 59668
rect 580276 59604 580277 59668
rect 580211 59603 580277 59604
rect 580214 48517 580274 59603
rect 580211 48516 580277 48517
rect 580211 48452 580212 48516
rect 580276 48452 580277 48516
rect 580211 48451 580277 48452
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16250 579218 16486 579454
rect 16250 578898 16486 579134
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16250 543218 16486 543454
rect 16250 542898 16486 543134
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16250 507218 16486 507454
rect 16250 506898 16486 507134
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16250 471218 16486 471454
rect 16250 470898 16486 471134
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16250 435218 16486 435454
rect 16250 434898 16486 435134
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16250 399218 16486 399454
rect 16250 398898 16486 399134
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16250 363218 16486 363454
rect 16250 362898 16486 363134
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16250 327218 16486 327454
rect 16250 326898 16486 327134
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16250 291218 16486 291454
rect 16250 290898 16486 291134
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16250 255218 16486 255454
rect 16250 254898 16486 255134
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16250 219218 16486 219454
rect 16250 218898 16486 219134
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16250 183218 16486 183454
rect 16250 182898 16486 183134
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16250 147218 16486 147454
rect 16250 146898 16486 147134
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16250 111218 16486 111454
rect 16250 110898 16486 111134
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16250 75218 16486 75454
rect 16250 74898 16486 75134
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16250 39218 16486 39454
rect 16250 38898 16486 39134
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 21370 582938 21606 583174
rect 21370 582618 21606 582854
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 26490 586658 26726 586894
rect 26490 586338 26726 586574
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 21370 546938 21606 547174
rect 21370 546618 21606 546854
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 36730 594098 36966 594334
rect 36730 593778 36966 594014
rect 31610 590378 31846 590614
rect 31610 590058 31846 590294
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 26490 550658 26726 550894
rect 26490 550338 26726 550574
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 21370 510938 21606 511174
rect 21370 510618 21606 510854
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 41850 597818 42086 598054
rect 41850 597498 42086 597734
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 36730 558098 36966 558334
rect 36730 557778 36966 558014
rect 31610 554378 31846 554614
rect 31610 554058 31846 554294
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 26490 514658 26726 514894
rect 26490 514338 26726 514574
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 21370 474938 21606 475174
rect 21370 474618 21606 474854
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 41850 561818 42086 562054
rect 41850 561498 42086 561734
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 36730 522098 36966 522334
rect 36730 521778 36966 522014
rect 31610 518378 31846 518614
rect 31610 518058 31846 518294
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 26490 478658 26726 478894
rect 26490 478338 26726 478574
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 21370 438938 21606 439174
rect 21370 438618 21606 438854
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 46970 579218 47206 579454
rect 46970 578898 47206 579134
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 41850 525818 42086 526054
rect 41850 525498 42086 525734
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 36730 486098 36966 486334
rect 36730 485778 36966 486014
rect 31610 482378 31846 482614
rect 31610 482058 31846 482294
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 26490 442658 26726 442894
rect 26490 442338 26726 442574
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 21370 402938 21606 403174
rect 21370 402618 21606 402854
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 52090 582938 52326 583174
rect 52090 582618 52326 582854
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 46970 543218 47206 543454
rect 46970 542898 47206 543134
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 41850 489818 42086 490054
rect 41850 489498 42086 489734
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 36730 450098 36966 450334
rect 36730 449778 36966 450014
rect 31610 446378 31846 446614
rect 31610 446058 31846 446294
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 26490 406658 26726 406894
rect 26490 406338 26726 406574
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 21370 366938 21606 367174
rect 21370 366618 21606 366854
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 52090 546938 52326 547174
rect 52090 546618 52326 546854
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 46970 507218 47206 507454
rect 46970 506898 47206 507134
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 41850 453818 42086 454054
rect 41850 453498 42086 453734
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 36730 414098 36966 414334
rect 36730 413778 36966 414014
rect 31610 410378 31846 410614
rect 31610 410058 31846 410294
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 26490 370658 26726 370894
rect 26490 370338 26726 370574
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 21370 330938 21606 331174
rect 21370 330618 21606 330854
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 52090 510938 52326 511174
rect 52090 510618 52326 510854
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 46970 471218 47206 471454
rect 46970 470898 47206 471134
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 41850 417818 42086 418054
rect 41850 417498 42086 417734
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 36730 378098 36966 378334
rect 36730 377778 36966 378014
rect 31610 374378 31846 374614
rect 31610 374058 31846 374294
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 26490 334658 26726 334894
rect 26490 334338 26726 334574
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 21370 294938 21606 295174
rect 21370 294618 21606 294854
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52090 474938 52326 475174
rect 52090 474618 52326 474854
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 46970 435218 47206 435454
rect 46970 434898 47206 435134
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 41850 381818 42086 382054
rect 41850 381498 42086 381734
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 36730 342098 36966 342334
rect 36730 341778 36966 342014
rect 31610 338378 31846 338614
rect 31610 338058 31846 338294
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 26490 298658 26726 298894
rect 26490 298338 26726 298574
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 21370 258938 21606 259174
rect 21370 258618 21606 258854
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52090 438938 52326 439174
rect 52090 438618 52326 438854
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 46970 399218 47206 399454
rect 46970 398898 47206 399134
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 41850 345818 42086 346054
rect 41850 345498 42086 345734
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 36730 306098 36966 306334
rect 36730 305778 36966 306014
rect 31610 302378 31846 302614
rect 31610 302058 31846 302294
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 26490 262658 26726 262894
rect 26490 262338 26726 262574
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 21370 222938 21606 223174
rect 21370 222618 21606 222854
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52090 402938 52326 403174
rect 52090 402618 52326 402854
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 46970 363218 47206 363454
rect 46970 362898 47206 363134
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 41850 309818 42086 310054
rect 41850 309498 42086 309734
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 36730 270098 36966 270334
rect 36730 269778 36966 270014
rect 31610 266378 31846 266614
rect 31610 266058 31846 266294
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 26490 226658 26726 226894
rect 26490 226338 26726 226574
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 21370 186938 21606 187174
rect 21370 186618 21606 186854
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52090 366938 52326 367174
rect 52090 366618 52326 366854
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 46970 327218 47206 327454
rect 46970 326898 47206 327134
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 41850 273818 42086 274054
rect 41850 273498 42086 273734
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 36730 234098 36966 234334
rect 36730 233778 36966 234014
rect 31610 230378 31846 230614
rect 31610 230058 31846 230294
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 26490 190658 26726 190894
rect 26490 190338 26726 190574
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 21370 150938 21606 151174
rect 21370 150618 21606 150854
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52090 330938 52326 331174
rect 52090 330618 52326 330854
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 46970 291218 47206 291454
rect 46970 290898 47206 291134
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 41850 237818 42086 238054
rect 41850 237498 42086 237734
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 36730 198098 36966 198334
rect 36730 197778 36966 198014
rect 31610 194378 31846 194614
rect 31610 194058 31846 194294
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 26490 154658 26726 154894
rect 26490 154338 26726 154574
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 21370 114938 21606 115174
rect 21370 114618 21606 114854
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 52090 294938 52326 295174
rect 52090 294618 52326 294854
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 46970 255218 47206 255454
rect 46970 254898 47206 255134
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 41850 201818 42086 202054
rect 41850 201498 42086 201734
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 36730 162098 36966 162334
rect 36730 161778 36966 162014
rect 31610 158378 31846 158614
rect 31610 158058 31846 158294
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 26490 118658 26726 118894
rect 26490 118338 26726 118574
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 21370 78938 21606 79174
rect 21370 78618 21606 78854
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 52090 258938 52326 259174
rect 52090 258618 52326 258854
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 46970 219218 47206 219454
rect 46970 218898 47206 219134
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 41850 165818 42086 166054
rect 41850 165498 42086 165734
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 36730 126098 36966 126334
rect 36730 125778 36966 126014
rect 31610 122378 31846 122614
rect 31610 122058 31846 122294
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 26490 82658 26726 82894
rect 26490 82338 26726 82574
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 21370 42938 21606 43174
rect 21370 42618 21606 42854
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52090 222938 52326 223174
rect 52090 222618 52326 222854
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 46970 183218 47206 183454
rect 46970 182898 47206 183134
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 41850 129818 42086 130054
rect 41850 129498 42086 129734
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 36730 90098 36966 90334
rect 36730 89778 36966 90014
rect 31610 86378 31846 86614
rect 31610 86058 31846 86294
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 26490 46658 26726 46894
rect 26490 46338 26726 46574
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 21370 6938 21606 7174
rect 21370 6618 21606 6854
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52090 186938 52326 187174
rect 52090 186618 52326 186854
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 46970 147218 47206 147454
rect 46970 146898 47206 147134
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 41850 93818 42086 94054
rect 41850 93498 42086 93734
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 36730 54098 36966 54334
rect 36730 53778 36966 54014
rect 31610 50378 31846 50614
rect 31610 50058 31846 50294
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 26490 10658 26726 10894
rect 26490 10338 26726 10574
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 52090 150938 52326 151174
rect 52090 150618 52326 150854
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 46970 111218 47206 111454
rect 46970 110898 47206 111134
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 41850 57818 42086 58054
rect 41850 57498 42086 57734
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 36730 18098 36966 18334
rect 36730 17778 36966 18014
rect 31610 14378 31846 14614
rect 31610 14058 31846 14294
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 52090 114938 52326 115174
rect 52090 114618 52326 114854
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 46970 75218 47206 75454
rect 46970 74898 47206 75134
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 41850 21818 42086 22054
rect 41850 21498 42086 21734
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 52090 78938 52326 79174
rect 52090 78618 52326 78854
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 46970 39218 47206 39454
rect 46970 38898 47206 39134
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52090 42938 52326 43174
rect 52090 42618 52326 42854
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52090 6938 52326 7174
rect 52090 6618 52326 6854
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 57210 586658 57446 586894
rect 57210 586338 57446 586574
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 63866 605258 64102 605494
rect 64186 605258 64422 605494
rect 63866 604938 64102 605174
rect 64186 604938 64422 605174
rect 62330 590378 62566 590614
rect 62330 590058 62566 590294
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 57210 550658 57446 550894
rect 57210 550338 57446 550574
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 72570 597818 72806 598054
rect 72570 597498 72806 597734
rect 67450 594098 67686 594334
rect 67450 593778 67686 594014
rect 63866 569258 64102 569494
rect 64186 569258 64422 569494
rect 63866 568938 64102 569174
rect 64186 568938 64422 569174
rect 62330 554378 62566 554614
rect 62330 554058 62566 554294
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 57210 514658 57446 514894
rect 57210 514338 57446 514574
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 72570 561818 72806 562054
rect 72570 561498 72806 561734
rect 67450 558098 67686 558334
rect 67450 557778 67686 558014
rect 63866 533258 64102 533494
rect 64186 533258 64422 533494
rect 63866 532938 64102 533174
rect 64186 532938 64422 533174
rect 62330 518378 62566 518614
rect 62330 518058 62566 518294
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 57210 478658 57446 478894
rect 57210 478338 57446 478574
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 77690 579218 77926 579454
rect 77690 578898 77926 579134
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 82810 582938 83046 583174
rect 82810 582618 83046 582854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 72570 525818 72806 526054
rect 72570 525498 72806 525734
rect 67450 522098 67686 522334
rect 67450 521778 67686 522014
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 62330 482378 62566 482614
rect 62330 482058 62566 482294
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 57210 442658 57446 442894
rect 57210 442338 57446 442574
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 77690 543218 77926 543454
rect 77690 542898 77926 543134
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 88706 630098 88942 630334
rect 89026 630098 89262 630334
rect 88706 629778 88942 630014
rect 89026 629778 89262 630014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 88706 594098 88942 594334
rect 89026 594098 89262 594334
rect 88706 593778 88942 594014
rect 89026 593778 89262 594014
rect 87930 586658 88166 586894
rect 87930 586338 88166 586574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 82810 546938 83046 547174
rect 82810 546618 83046 546854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 72570 489818 72806 490054
rect 72570 489498 72806 489734
rect 67450 486098 67686 486334
rect 67450 485778 67686 486014
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 62330 446378 62566 446614
rect 62330 446058 62566 446294
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 57210 406658 57446 406894
rect 57210 406338 57446 406574
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 77690 507218 77926 507454
rect 77690 506898 77926 507134
rect 96146 601538 96382 601774
rect 96466 601538 96702 601774
rect 96146 601218 96382 601454
rect 96466 601218 96702 601454
rect 93050 590378 93286 590614
rect 93050 590058 93286 590294
rect 88706 558098 88942 558334
rect 89026 558098 89262 558334
rect 88706 557778 88942 558014
rect 89026 557778 89262 558014
rect 87930 550658 88166 550894
rect 87930 550338 88166 550574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 82810 510938 83046 511174
rect 82810 510618 83046 510854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 72570 453818 72806 454054
rect 72570 453498 72806 453734
rect 67450 450098 67686 450334
rect 67450 449778 67686 450014
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 62330 410378 62566 410614
rect 62330 410058 62566 410294
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 57210 370658 57446 370894
rect 57210 370338 57446 370574
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 77690 471218 77926 471454
rect 77690 470898 77926 471134
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 99866 605258 100102 605494
rect 100186 605258 100422 605494
rect 99866 604938 100102 605174
rect 100186 604938 100422 605174
rect 98170 594098 98406 594334
rect 98170 593778 98406 594014
rect 96146 565538 96382 565774
rect 96466 565538 96702 565774
rect 96146 565218 96382 565454
rect 96466 565218 96702 565454
rect 93050 554378 93286 554614
rect 93050 554058 93286 554294
rect 88706 522098 88942 522334
rect 89026 522098 89262 522334
rect 88706 521778 88942 522014
rect 89026 521778 89262 522014
rect 87930 514658 88166 514894
rect 87930 514338 88166 514574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 82810 474938 83046 475174
rect 82810 474618 83046 474854
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 72570 417818 72806 418054
rect 72570 417498 72806 417734
rect 67450 414098 67686 414334
rect 67450 413778 67686 414014
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 62330 374378 62566 374614
rect 62330 374058 62566 374294
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 57210 334658 57446 334894
rect 57210 334338 57446 334574
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 77690 435218 77926 435454
rect 77690 434898 77926 435134
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 103290 597818 103526 598054
rect 103290 597498 103526 597734
rect 108410 579218 108646 579454
rect 108410 578898 108646 579134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 124706 630098 124942 630334
rect 125026 630098 125262 630334
rect 124706 629778 124942 630014
rect 125026 629778 125262 630014
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 132146 601538 132382 601774
rect 132466 601538 132702 601774
rect 132146 601218 132382 601454
rect 132466 601218 132702 601454
rect 124706 594098 124942 594334
rect 125026 594098 125262 594334
rect 124706 593778 124942 594014
rect 125026 593778 125262 594014
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 113530 582938 113766 583174
rect 113530 582618 113766 582854
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 99866 569258 100102 569494
rect 100186 569258 100422 569494
rect 99866 568938 100102 569174
rect 100186 568938 100422 569174
rect 98170 558098 98406 558334
rect 98170 557778 98406 558014
rect 96146 529538 96382 529774
rect 96466 529538 96702 529774
rect 96146 529218 96382 529454
rect 96466 529218 96702 529454
rect 93050 518378 93286 518614
rect 93050 518058 93286 518294
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 87930 478658 88166 478894
rect 87930 478338 88166 478574
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 82810 438938 83046 439174
rect 82810 438618 83046 438854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 72570 381818 72806 382054
rect 72570 381498 72806 381734
rect 67450 378098 67686 378334
rect 67450 377778 67686 378014
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 62330 338378 62566 338614
rect 62330 338058 62566 338294
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 57210 298658 57446 298894
rect 57210 298338 57446 298574
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 77690 399218 77926 399454
rect 77690 398898 77926 399134
rect 103290 561818 103526 562054
rect 103290 561498 103526 561734
rect 108410 543218 108646 543454
rect 108410 542898 108646 543134
rect 118650 586658 118886 586894
rect 118650 586338 118886 586574
rect 123770 590378 124006 590614
rect 123770 590058 124006 590294
rect 128890 594098 129126 594334
rect 128890 593778 129126 594014
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 135866 605258 136102 605494
rect 136186 605258 136422 605494
rect 135866 604938 136102 605174
rect 136186 604938 136422 605174
rect 134010 597818 134246 598054
rect 134010 597498 134246 597734
rect 132146 565538 132382 565774
rect 132466 565538 132702 565774
rect 132146 565218 132382 565454
rect 132466 565218 132702 565454
rect 124706 558098 124942 558334
rect 125026 558098 125262 558334
rect 124706 557778 124942 558014
rect 125026 557778 125262 558014
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 113530 546938 113766 547174
rect 113530 546618 113766 546854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 99866 533258 100102 533494
rect 100186 533258 100422 533494
rect 99866 532938 100102 533174
rect 100186 532938 100422 533174
rect 98170 522098 98406 522334
rect 98170 521778 98406 522014
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 93050 482378 93286 482614
rect 93050 482058 93286 482294
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 87930 442658 88166 442894
rect 87930 442338 88166 442574
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 82810 402938 83046 403174
rect 82810 402618 83046 402854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 72570 345818 72806 346054
rect 72570 345498 72806 345734
rect 67450 342098 67686 342334
rect 67450 341778 67686 342014
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 62330 302378 62566 302614
rect 62330 302058 62566 302294
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 57210 262658 57446 262894
rect 57210 262338 57446 262574
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 77690 363218 77926 363454
rect 77690 362898 77926 363134
rect 103290 525818 103526 526054
rect 103290 525498 103526 525734
rect 108410 507218 108646 507454
rect 108410 506898 108646 507134
rect 118650 550658 118886 550894
rect 118650 550338 118886 550574
rect 123770 554378 124006 554614
rect 123770 554058 124006 554294
rect 128890 558098 129126 558334
rect 128890 557778 129126 558014
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 144250 582938 144486 583174
rect 144250 582618 144486 582854
rect 139130 579218 139366 579454
rect 139130 578898 139366 579134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 149370 586658 149606 586894
rect 149370 586338 149606 586574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 154490 590378 154726 590614
rect 154490 590058 154726 590294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 159610 594098 159846 594334
rect 159610 593778 159846 594014
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 164730 597818 164966 598054
rect 164730 597498 164966 597734
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 135866 569258 136102 569494
rect 136186 569258 136422 569494
rect 135866 568938 136102 569174
rect 136186 568938 136422 569174
rect 134010 561818 134246 562054
rect 134010 561498 134246 561734
rect 132146 529538 132382 529774
rect 132466 529538 132702 529774
rect 132146 529218 132382 529454
rect 132466 529218 132702 529454
rect 124706 522098 124942 522334
rect 125026 522098 125262 522334
rect 124706 521778 124942 522014
rect 125026 521778 125262 522014
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 113530 510938 113766 511174
rect 113530 510618 113766 510854
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 98170 486098 98406 486334
rect 98170 485778 98406 486014
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 93050 446378 93286 446614
rect 93050 446058 93286 446294
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 87930 406658 88166 406894
rect 87930 406338 88166 406574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 82810 366938 83046 367174
rect 82810 366618 83046 366854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 72570 309818 72806 310054
rect 72570 309498 72806 309734
rect 67450 306098 67686 306334
rect 67450 305778 67686 306014
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 62330 266378 62566 266614
rect 62330 266058 62566 266294
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 57210 226658 57446 226894
rect 57210 226338 57446 226574
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 77690 327218 77926 327454
rect 77690 326898 77926 327134
rect 103290 489818 103526 490054
rect 103290 489498 103526 489734
rect 108410 471218 108646 471454
rect 108410 470898 108646 471134
rect 118650 514658 118886 514894
rect 118650 514338 118886 514574
rect 123770 518378 124006 518614
rect 123770 518058 124006 518294
rect 128890 522098 129126 522334
rect 128890 521778 129126 522014
rect 144250 546938 144486 547174
rect 144250 546618 144486 546854
rect 139130 543218 139366 543454
rect 139130 542898 139366 543134
rect 149370 550658 149606 550894
rect 149370 550338 149606 550574
rect 154490 554378 154726 554614
rect 154490 554058 154726 554294
rect 159610 558098 159846 558334
rect 159610 557778 159846 558014
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 169850 579218 170086 579454
rect 169850 578898 170086 579134
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 164730 561818 164966 562054
rect 164730 561498 164966 561734
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 135866 533258 136102 533494
rect 136186 533258 136422 533494
rect 135866 532938 136102 533174
rect 136186 532938 136422 533174
rect 134010 525818 134246 526054
rect 134010 525498 134246 525734
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113530 474938 113766 475174
rect 113530 474618 113766 474854
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 98170 450098 98406 450334
rect 98170 449778 98406 450014
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 93050 410378 93286 410614
rect 93050 410058 93286 410294
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 87930 370658 88166 370894
rect 87930 370338 88166 370574
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 82810 330938 83046 331174
rect 82810 330618 83046 330854
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 72570 273818 72806 274054
rect 72570 273498 72806 273734
rect 67450 270098 67686 270334
rect 67450 269778 67686 270014
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 62330 230378 62566 230614
rect 62330 230058 62566 230294
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 57210 190658 57446 190894
rect 57210 190338 57446 190574
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 77690 291218 77926 291454
rect 77690 290898 77926 291134
rect 103290 453818 103526 454054
rect 103290 453498 103526 453734
rect 108410 435218 108646 435454
rect 108410 434898 108646 435134
rect 118650 478658 118886 478894
rect 118650 478338 118886 478574
rect 123770 482378 124006 482614
rect 123770 482058 124006 482294
rect 128890 486098 129126 486334
rect 128890 485778 129126 486014
rect 144250 510938 144486 511174
rect 144250 510618 144486 510854
rect 139130 507218 139366 507454
rect 139130 506898 139366 507134
rect 149370 514658 149606 514894
rect 149370 514338 149606 514574
rect 154490 518378 154726 518614
rect 154490 518058 154726 518294
rect 159610 522098 159846 522334
rect 159610 521778 159846 522014
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 180090 586658 180326 586894
rect 180090 586338 180326 586574
rect 174970 582938 175206 583174
rect 174970 582618 175206 582854
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 169850 543218 170086 543454
rect 169850 542898 170086 543134
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 164730 525818 164966 526054
rect 164730 525498 164966 525734
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 134010 489818 134246 490054
rect 134010 489498 134246 489734
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 113530 438938 113766 439174
rect 113530 438618 113766 438854
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 98170 414098 98406 414334
rect 98170 413778 98406 414014
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 93050 374378 93286 374614
rect 93050 374058 93286 374294
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 87930 334658 88166 334894
rect 87930 334338 88166 334574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 82810 294938 83046 295174
rect 82810 294618 83046 294854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 72570 237818 72806 238054
rect 72570 237498 72806 237734
rect 67450 234098 67686 234334
rect 67450 233778 67686 234014
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 62330 194378 62566 194614
rect 62330 194058 62566 194294
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 57210 154658 57446 154894
rect 57210 154338 57446 154574
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 77690 255218 77926 255454
rect 77690 254898 77926 255134
rect 103290 417818 103526 418054
rect 103290 417498 103526 417734
rect 108410 399218 108646 399454
rect 108410 398898 108646 399134
rect 118650 442658 118886 442894
rect 118650 442338 118886 442574
rect 123770 446378 124006 446614
rect 123770 446058 124006 446294
rect 128890 450098 129126 450334
rect 128890 449778 129126 450014
rect 144250 474938 144486 475174
rect 144250 474618 144486 474854
rect 139130 471218 139366 471454
rect 139130 470898 139366 471134
rect 149370 478658 149606 478894
rect 149370 478338 149606 478574
rect 154490 482378 154726 482614
rect 154490 482058 154726 482294
rect 159610 486098 159846 486334
rect 159610 485778 159846 486014
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 185210 590378 185446 590614
rect 185210 590058 185446 590294
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 180090 550658 180326 550894
rect 180090 550338 180326 550574
rect 174970 546938 175206 547174
rect 174970 546618 175206 546854
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 169850 507218 170086 507454
rect 169850 506898 170086 507134
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 164730 489818 164966 490054
rect 164730 489498 164966 489734
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 134010 453818 134246 454054
rect 134010 453498 134246 453734
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 113530 402938 113766 403174
rect 113530 402618 113766 402854
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 98170 378098 98406 378334
rect 98170 377778 98406 378014
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 93050 338378 93286 338614
rect 93050 338058 93286 338294
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 87930 298658 88166 298894
rect 87930 298338 88166 298574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 82810 258938 83046 259174
rect 82810 258618 83046 258854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 72570 201818 72806 202054
rect 72570 201498 72806 201734
rect 67450 198098 67686 198334
rect 67450 197778 67686 198014
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 62330 158378 62566 158614
rect 62330 158058 62566 158294
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 57210 118658 57446 118894
rect 57210 118338 57446 118574
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 77690 219218 77926 219454
rect 77690 218898 77926 219134
rect 103290 381818 103526 382054
rect 103290 381498 103526 381734
rect 108410 363218 108646 363454
rect 108410 362898 108646 363134
rect 118650 406658 118886 406894
rect 118650 406338 118886 406574
rect 123770 410378 124006 410614
rect 123770 410058 124006 410294
rect 128890 414098 129126 414334
rect 128890 413778 129126 414014
rect 144250 438938 144486 439174
rect 144250 438618 144486 438854
rect 139130 435218 139366 435454
rect 139130 434898 139366 435134
rect 149370 442658 149606 442894
rect 149370 442338 149606 442574
rect 154490 446378 154726 446614
rect 154490 446058 154726 446294
rect 159610 450098 159846 450334
rect 159610 449778 159846 450014
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 190330 594098 190566 594334
rect 190330 593778 190566 594014
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 185210 554378 185446 554614
rect 185210 554058 185446 554294
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 180090 514658 180326 514894
rect 180090 514338 180326 514574
rect 174970 510938 175206 511174
rect 174970 510618 175206 510854
rect 171866 497258 172102 497494
rect 172186 497258 172422 497494
rect 171866 496938 172102 497174
rect 172186 496938 172422 497174
rect 169850 471218 170086 471454
rect 169850 470898 170086 471134
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 164730 453818 164966 454054
rect 164730 453498 164966 453734
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 134010 417818 134246 418054
rect 134010 417498 134246 417734
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 113530 366938 113766 367174
rect 113530 366618 113766 366854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 98170 342098 98406 342334
rect 98170 341778 98406 342014
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 93050 302378 93286 302614
rect 93050 302058 93286 302294
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 87930 262658 88166 262894
rect 87930 262338 88166 262574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 82810 222938 83046 223174
rect 82810 222618 83046 222854
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 72570 165818 72806 166054
rect 72570 165498 72806 165734
rect 67450 162098 67686 162334
rect 67450 161778 67686 162014
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 62330 122378 62566 122614
rect 62330 122058 62566 122294
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 57210 82658 57446 82894
rect 57210 82338 57446 82574
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 77690 183218 77926 183454
rect 77690 182898 77926 183134
rect 103290 345818 103526 346054
rect 103290 345498 103526 345734
rect 108410 327218 108646 327454
rect 108410 326898 108646 327134
rect 118650 370658 118886 370894
rect 118650 370338 118886 370574
rect 123770 374378 124006 374614
rect 123770 374058 124006 374294
rect 128890 378098 129126 378334
rect 128890 377778 129126 378014
rect 144250 402938 144486 403174
rect 144250 402618 144486 402854
rect 139130 399218 139366 399454
rect 139130 398898 139366 399134
rect 149370 406658 149606 406894
rect 149370 406338 149606 406574
rect 154490 410378 154726 410614
rect 154490 410058 154726 410294
rect 159610 414098 159846 414334
rect 159610 413778 159846 414014
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 195450 597818 195686 598054
rect 195450 597498 195686 597734
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 190330 558098 190566 558334
rect 190330 557778 190566 558014
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 185210 518378 185446 518614
rect 185210 518058 185446 518294
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 180090 478658 180326 478894
rect 180090 478338 180326 478574
rect 174970 474938 175206 475174
rect 174970 474618 175206 474854
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 169850 435218 170086 435454
rect 169850 434898 170086 435134
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 164730 417818 164966 418054
rect 164730 417498 164966 417734
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 134010 381818 134246 382054
rect 134010 381498 134246 381734
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 113530 330938 113766 331174
rect 113530 330618 113766 330854
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 98170 306098 98406 306334
rect 98170 305778 98406 306014
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 93050 266378 93286 266614
rect 93050 266058 93286 266294
rect 88706 234098 88942 234334
rect 89026 234098 89262 234334
rect 88706 233778 88942 234014
rect 89026 233778 89262 234014
rect 87930 226658 88166 226894
rect 87930 226338 88166 226574
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 82810 186938 83046 187174
rect 82810 186618 83046 186854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 72570 129818 72806 130054
rect 72570 129498 72806 129734
rect 67450 126098 67686 126334
rect 67450 125778 67686 126014
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 62330 86378 62566 86614
rect 62330 86058 62566 86294
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 57210 46658 57446 46894
rect 57210 46338 57446 46574
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 77690 147218 77926 147454
rect 77690 146898 77926 147134
rect 103290 309818 103526 310054
rect 103290 309498 103526 309734
rect 108410 291218 108646 291454
rect 108410 290898 108646 291134
rect 118650 334658 118886 334894
rect 118650 334338 118886 334574
rect 123770 338378 124006 338614
rect 123770 338058 124006 338294
rect 128890 342098 129126 342334
rect 128890 341778 129126 342014
rect 144250 366938 144486 367174
rect 144250 366618 144486 366854
rect 139130 363218 139366 363454
rect 139130 362898 139366 363134
rect 149370 370658 149606 370894
rect 149370 370338 149606 370574
rect 154490 374378 154726 374614
rect 154490 374058 154726 374294
rect 159610 378098 159846 378334
rect 159610 377778 159846 378014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 195450 561818 195686 562054
rect 195450 561498 195686 561734
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 190330 522098 190566 522334
rect 190330 521778 190566 522014
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 185210 482378 185446 482614
rect 185210 482058 185446 482294
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 180090 442658 180326 442894
rect 180090 442338 180326 442574
rect 174970 438938 175206 439174
rect 174970 438618 175206 438854
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 169850 399218 170086 399454
rect 169850 398898 170086 399134
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 164730 381818 164966 382054
rect 164730 381498 164966 381734
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 134010 345818 134246 346054
rect 134010 345498 134246 345734
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 113530 294938 113766 295174
rect 113530 294618 113766 294854
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 99866 281258 100102 281494
rect 100186 281258 100422 281494
rect 99866 280938 100102 281174
rect 100186 280938 100422 281174
rect 98170 270098 98406 270334
rect 98170 269778 98406 270014
rect 96146 241538 96382 241774
rect 96466 241538 96702 241774
rect 96146 241218 96382 241454
rect 96466 241218 96702 241454
rect 93050 230378 93286 230614
rect 93050 230058 93286 230294
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 87930 190658 88166 190894
rect 87930 190338 88166 190574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 82810 150938 83046 151174
rect 82810 150618 83046 150854
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 72570 93818 72806 94054
rect 72570 93498 72806 93734
rect 67450 90098 67686 90334
rect 67450 89778 67686 90014
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 62330 50378 62566 50614
rect 62330 50058 62566 50294
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 57210 10658 57446 10894
rect 57210 10338 57446 10574
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 77690 111218 77926 111454
rect 77690 110898 77926 111134
rect 103290 273818 103526 274054
rect 103290 273498 103526 273734
rect 108410 255218 108646 255454
rect 108410 254898 108646 255134
rect 118650 298658 118886 298894
rect 118650 298338 118886 298574
rect 123770 302378 124006 302614
rect 123770 302058 124006 302294
rect 128890 306098 129126 306334
rect 128890 305778 129126 306014
rect 144250 330938 144486 331174
rect 144250 330618 144486 330854
rect 139130 327218 139366 327454
rect 139130 326898 139366 327134
rect 149370 334658 149606 334894
rect 149370 334338 149606 334574
rect 154490 338378 154726 338614
rect 154490 338058 154726 338294
rect 159610 342098 159846 342334
rect 159610 341778 159846 342014
rect 204146 601538 204382 601774
rect 204466 601538 204702 601774
rect 204146 601218 204382 601454
rect 204466 601218 204702 601454
rect 200570 579218 200806 579454
rect 200570 578898 200806 579134
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 195450 525818 195686 526054
rect 195450 525498 195686 525734
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 190330 486098 190566 486334
rect 190330 485778 190566 486014
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 185210 446378 185446 446614
rect 185210 446058 185446 446294
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 180090 406658 180326 406894
rect 180090 406338 180326 406574
rect 174970 402938 175206 403174
rect 174970 402618 175206 402854
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 169850 363218 170086 363454
rect 169850 362898 170086 363134
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 164730 345818 164966 346054
rect 164730 345498 164966 345734
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 134010 309818 134246 310054
rect 134010 309498 134246 309734
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 113530 258938 113766 259174
rect 113530 258618 113766 258854
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 99866 245258 100102 245494
rect 100186 245258 100422 245494
rect 99866 244938 100102 245174
rect 100186 244938 100422 245174
rect 98170 234098 98406 234334
rect 98170 233778 98406 234014
rect 96146 205538 96382 205774
rect 96466 205538 96702 205774
rect 96146 205218 96382 205454
rect 96466 205218 96702 205454
rect 93050 194378 93286 194614
rect 93050 194058 93286 194294
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 87930 154658 88166 154894
rect 87930 154338 88166 154574
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 82810 114938 83046 115174
rect 82810 114618 83046 114854
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 72570 57818 72806 58054
rect 72570 57498 72806 57734
rect 67450 54098 67686 54334
rect 67450 53778 67686 54014
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 62330 14378 62566 14614
rect 62330 14058 62566 14294
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 77690 75218 77926 75454
rect 77690 74898 77926 75134
rect 103290 237818 103526 238054
rect 103290 237498 103526 237734
rect 108410 219218 108646 219454
rect 108410 218898 108646 219134
rect 118650 262658 118886 262894
rect 118650 262338 118886 262574
rect 123770 266378 124006 266614
rect 123770 266058 124006 266294
rect 128890 270098 129126 270334
rect 128890 269778 129126 270014
rect 144250 294938 144486 295174
rect 144250 294618 144486 294854
rect 139130 291218 139366 291454
rect 139130 290898 139366 291134
rect 149370 298658 149606 298894
rect 149370 298338 149606 298574
rect 154490 302378 154726 302614
rect 154490 302058 154726 302294
rect 159610 306098 159846 306334
rect 159610 305778 159846 306014
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 205690 582938 205926 583174
rect 205690 582618 205926 582854
rect 204146 565538 204382 565774
rect 204466 565538 204702 565774
rect 204146 565218 204382 565454
rect 204466 565218 204702 565454
rect 200570 543218 200806 543454
rect 200570 542898 200806 543134
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 195450 489818 195686 490054
rect 195450 489498 195686 489734
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 190330 450098 190566 450334
rect 190330 449778 190566 450014
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 185210 410378 185446 410614
rect 185210 410058 185446 410294
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 180090 370658 180326 370894
rect 180090 370338 180326 370574
rect 174970 366938 175206 367174
rect 174970 366618 175206 366854
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 169850 327218 170086 327454
rect 169850 326898 170086 327134
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 164730 309818 164966 310054
rect 164730 309498 164966 309734
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 134010 273818 134246 274054
rect 134010 273498 134246 273734
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 113530 222938 113766 223174
rect 113530 222618 113766 222854
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 99866 209258 100102 209494
rect 100186 209258 100422 209494
rect 99866 208938 100102 209174
rect 100186 208938 100422 209174
rect 98170 198098 98406 198334
rect 98170 197778 98406 198014
rect 96146 169538 96382 169774
rect 96466 169538 96702 169774
rect 96146 169218 96382 169454
rect 96466 169218 96702 169454
rect 93050 158378 93286 158614
rect 93050 158058 93286 158294
rect 88706 126098 88942 126334
rect 89026 126098 89262 126334
rect 88706 125778 88942 126014
rect 89026 125778 89262 126014
rect 87930 118658 88166 118894
rect 87930 118338 88166 118574
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 82810 78938 83046 79174
rect 82810 78618 83046 78854
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 72570 21818 72806 22054
rect 72570 21498 72806 21734
rect 67450 18098 67686 18334
rect 67450 17778 67686 18014
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 77690 39218 77926 39454
rect 77690 38898 77926 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 103290 201818 103526 202054
rect 103290 201498 103526 201734
rect 108410 183218 108646 183454
rect 108410 182898 108646 183134
rect 118650 226658 118886 226894
rect 118650 226338 118886 226574
rect 123770 230378 124006 230614
rect 123770 230058 124006 230294
rect 128890 234098 129126 234334
rect 128890 233778 129126 234014
rect 144250 258938 144486 259174
rect 144250 258618 144486 258854
rect 139130 255218 139366 255454
rect 139130 254898 139366 255134
rect 149370 262658 149606 262894
rect 149370 262338 149606 262574
rect 154490 266378 154726 266614
rect 154490 266058 154726 266294
rect 159610 270098 159846 270334
rect 159610 269778 159846 270014
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 215930 590378 216166 590614
rect 215930 590058 216166 590294
rect 210810 586658 211046 586894
rect 210810 586338 211046 586574
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 205690 546938 205926 547174
rect 205690 546618 205926 546854
rect 204146 529538 204382 529774
rect 204466 529538 204702 529774
rect 204146 529218 204382 529454
rect 204466 529218 204702 529454
rect 200570 507218 200806 507454
rect 200570 506898 200806 507134
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 195450 453818 195686 454054
rect 195450 453498 195686 453734
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 190330 414098 190566 414334
rect 190330 413778 190566 414014
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 185210 374378 185446 374614
rect 185210 374058 185446 374294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 180090 334658 180326 334894
rect 180090 334338 180326 334574
rect 174970 330938 175206 331174
rect 174970 330618 175206 330854
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 169850 291218 170086 291454
rect 169850 290898 170086 291134
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 164730 273818 164966 274054
rect 164730 273498 164966 273734
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 134010 237818 134246 238054
rect 134010 237498 134246 237734
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 113530 186938 113766 187174
rect 113530 186618 113766 186854
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 99866 173258 100102 173494
rect 100186 173258 100422 173494
rect 99866 172938 100102 173174
rect 100186 172938 100422 173174
rect 98170 162098 98406 162334
rect 98170 161778 98406 162014
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 93050 122378 93286 122614
rect 93050 122058 93286 122294
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 87930 82658 88166 82894
rect 87930 82338 88166 82574
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 82810 42938 83046 43174
rect 82810 42618 83046 42854
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 103290 165818 103526 166054
rect 103290 165498 103526 165734
rect 108410 147218 108646 147454
rect 108410 146898 108646 147134
rect 118650 190658 118886 190894
rect 118650 190338 118886 190574
rect 123770 194378 124006 194614
rect 123770 194058 124006 194294
rect 128890 198098 129126 198334
rect 128890 197778 129126 198014
rect 144250 222938 144486 223174
rect 144250 222618 144486 222854
rect 139130 219218 139366 219454
rect 139130 218898 139366 219134
rect 149370 226658 149606 226894
rect 149370 226338 149606 226574
rect 154490 230378 154726 230614
rect 154490 230058 154726 230294
rect 159610 234098 159846 234334
rect 159610 233778 159846 234014
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221050 594098 221286 594334
rect 221050 593778 221286 594014
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 215930 554378 216166 554614
rect 215930 554058 216166 554294
rect 210810 550658 211046 550894
rect 210810 550338 211046 550574
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 205690 510938 205926 511174
rect 205690 510618 205926 510854
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 200570 471218 200806 471454
rect 200570 470898 200806 471134
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 195450 417818 195686 418054
rect 195450 417498 195686 417734
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 190330 378098 190566 378334
rect 190330 377778 190566 378014
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 185210 338378 185446 338614
rect 185210 338058 185446 338294
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 180090 298658 180326 298894
rect 180090 298338 180326 298574
rect 174970 294938 175206 295174
rect 174970 294618 175206 294854
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 169850 255218 170086 255454
rect 169850 254898 170086 255134
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 164730 237818 164966 238054
rect 164730 237498 164966 237734
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 134010 201818 134246 202054
rect 134010 201498 134246 201734
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 113530 150938 113766 151174
rect 113530 150618 113766 150854
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 99866 137258 100102 137494
rect 100186 137258 100422 137494
rect 99866 136938 100102 137174
rect 100186 136938 100422 137174
rect 98170 126098 98406 126334
rect 98170 125778 98406 126014
rect 96146 97538 96382 97774
rect 96466 97538 96702 97774
rect 96146 97218 96382 97454
rect 96466 97218 96702 97454
rect 93050 86378 93286 86614
rect 93050 86058 93286 86294
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 87930 46658 88166 46894
rect 87930 46338 88166 46574
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 82810 6938 83046 7174
rect 82810 6618 83046 6854
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 103290 129818 103526 130054
rect 103290 129498 103526 129734
rect 108410 111218 108646 111454
rect 108410 110898 108646 111134
rect 118650 154658 118886 154894
rect 118650 154338 118886 154574
rect 123770 158378 124006 158614
rect 123770 158058 124006 158294
rect 128890 162098 129126 162334
rect 128890 161778 129126 162014
rect 144250 186938 144486 187174
rect 144250 186618 144486 186854
rect 139130 183218 139366 183454
rect 139130 182898 139366 183134
rect 149370 190658 149606 190894
rect 149370 190338 149606 190574
rect 154490 194378 154726 194614
rect 154490 194058 154726 194294
rect 159610 198098 159846 198334
rect 159610 197778 159846 198014
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221050 558098 221286 558334
rect 221050 557778 221286 558014
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 215930 518378 216166 518614
rect 215930 518058 216166 518294
rect 210810 514658 211046 514894
rect 210810 514338 211046 514574
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 205690 474938 205926 475174
rect 205690 474618 205926 474854
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 200570 435218 200806 435454
rect 200570 434898 200806 435134
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 195450 381818 195686 382054
rect 195450 381498 195686 381734
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 190330 342098 190566 342334
rect 190330 341778 190566 342014
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 185210 302378 185446 302614
rect 185210 302058 185446 302294
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 180090 262658 180326 262894
rect 180090 262338 180326 262574
rect 174970 258938 175206 259174
rect 174970 258618 175206 258854
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 169850 219218 170086 219454
rect 169850 218898 170086 219134
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 164730 201818 164966 202054
rect 164730 201498 164966 201734
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 134010 165818 134246 166054
rect 134010 165498 134246 165734
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 113530 114938 113766 115174
rect 113530 114618 113766 114854
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 99866 101258 100102 101494
rect 100186 101258 100422 101494
rect 99866 100938 100102 101174
rect 100186 100938 100422 101174
rect 98170 90098 98406 90334
rect 98170 89778 98406 90014
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 93050 50378 93286 50614
rect 93050 50058 93286 50294
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 87930 10658 88166 10894
rect 87930 10338 88166 10574
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 103290 93818 103526 94054
rect 103290 93498 103526 93734
rect 108410 75218 108646 75454
rect 108410 74898 108646 75134
rect 118650 118658 118886 118894
rect 118650 118338 118886 118574
rect 123770 122378 124006 122614
rect 123770 122058 124006 122294
rect 128890 126098 129126 126334
rect 128890 125778 129126 126014
rect 144250 150938 144486 151174
rect 144250 150618 144486 150854
rect 139130 147218 139366 147454
rect 139130 146898 139366 147134
rect 149370 154658 149606 154894
rect 149370 154338 149606 154574
rect 154490 158378 154726 158614
rect 154490 158058 154726 158294
rect 159610 162098 159846 162334
rect 159610 161778 159846 162014
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221050 522098 221286 522334
rect 221050 521778 221286 522014
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 215930 482378 216166 482614
rect 215930 482058 216166 482294
rect 210810 478658 211046 478894
rect 210810 478338 211046 478574
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 205690 438938 205926 439174
rect 205690 438618 205926 438854
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 200570 399218 200806 399454
rect 200570 398898 200806 399134
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 195450 345818 195686 346054
rect 195450 345498 195686 345734
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 190330 306098 190566 306334
rect 190330 305778 190566 306014
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 185210 266378 185446 266614
rect 185210 266058 185446 266294
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 180090 226658 180326 226894
rect 180090 226338 180326 226574
rect 174970 222938 175206 223174
rect 174970 222618 175206 222854
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 169850 183218 170086 183454
rect 169850 182898 170086 183134
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 164730 165818 164966 166054
rect 164730 165498 164966 165734
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 134010 129818 134246 130054
rect 134010 129498 134246 129734
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 113530 78938 113766 79174
rect 113530 78618 113766 78854
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 98170 54098 98406 54334
rect 98170 53778 98406 54014
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 93050 14378 93286 14614
rect 93050 14058 93286 14294
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 103290 57818 103526 58054
rect 103290 57498 103526 57734
rect 108410 39218 108646 39454
rect 108410 38898 108646 39134
rect 118650 82658 118886 82894
rect 118650 82338 118886 82574
rect 123770 86378 124006 86614
rect 123770 86058 124006 86294
rect 128890 90098 129126 90334
rect 128890 89778 129126 90014
rect 144250 114938 144486 115174
rect 144250 114618 144486 114854
rect 139130 111218 139366 111454
rect 139130 110898 139366 111134
rect 149370 118658 149606 118894
rect 149370 118338 149606 118574
rect 154490 122378 154726 122614
rect 154490 122058 154726 122294
rect 159610 126098 159846 126334
rect 159610 125778 159846 126014
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221050 486098 221286 486334
rect 221050 485778 221286 486014
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 215930 446378 216166 446614
rect 215930 446058 216166 446294
rect 210810 442658 211046 442894
rect 210810 442338 211046 442574
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 205690 402938 205926 403174
rect 205690 402618 205926 402854
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 200570 363218 200806 363454
rect 200570 362898 200806 363134
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 195450 309818 195686 310054
rect 195450 309498 195686 309734
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 190330 270098 190566 270334
rect 190330 269778 190566 270014
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 185210 230378 185446 230614
rect 185210 230058 185446 230294
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 180090 190658 180326 190894
rect 180090 190338 180326 190574
rect 174970 186938 175206 187174
rect 174970 186618 175206 186854
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 169850 147218 170086 147454
rect 169850 146898 170086 147134
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 164730 129818 164966 130054
rect 164730 129498 164966 129734
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 134010 93818 134246 94054
rect 134010 93498 134246 93734
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 113530 42938 113766 43174
rect 113530 42618 113766 42854
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 98170 18098 98406 18334
rect 98170 17778 98406 18014
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 103290 21818 103526 22054
rect 103290 21498 103526 21734
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 118650 46658 118886 46894
rect 118650 46338 118886 46574
rect 123770 50378 124006 50614
rect 123770 50058 124006 50294
rect 128890 54098 129126 54334
rect 128890 53778 129126 54014
rect 144250 78938 144486 79174
rect 144250 78618 144486 78854
rect 139130 75218 139366 75454
rect 139130 74898 139366 75134
rect 149370 82658 149606 82894
rect 149370 82338 149606 82574
rect 154490 86378 154726 86614
rect 154490 86058 154726 86294
rect 159610 90098 159846 90334
rect 159610 89778 159846 90014
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221050 450098 221286 450334
rect 221050 449778 221286 450014
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 215930 410378 216166 410614
rect 215930 410058 216166 410294
rect 210810 406658 211046 406894
rect 210810 406338 211046 406574
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 205690 366938 205926 367174
rect 205690 366618 205926 366854
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 200570 327218 200806 327454
rect 200570 326898 200806 327134
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 195450 273818 195686 274054
rect 195450 273498 195686 273734
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 190330 234098 190566 234334
rect 190330 233778 190566 234014
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 185210 194378 185446 194614
rect 185210 194058 185446 194294
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 180090 154658 180326 154894
rect 180090 154338 180326 154574
rect 174970 150938 175206 151174
rect 174970 150618 175206 150854
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 169850 111218 170086 111454
rect 169850 110898 170086 111134
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 164730 93818 164966 94054
rect 164730 93498 164966 93734
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 134010 57818 134246 58054
rect 134010 57498 134246 57734
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 113530 6938 113766 7174
rect 113530 6618 113766 6854
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 118650 10658 118886 10894
rect 118650 10338 118886 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 123770 14378 124006 14614
rect 123770 14058 124006 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 128890 18098 129126 18334
rect 128890 17778 129126 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 144250 42938 144486 43174
rect 144250 42618 144486 42854
rect 139130 39218 139366 39454
rect 139130 38898 139366 39134
rect 149370 46658 149606 46894
rect 149370 46338 149606 46574
rect 154490 50378 154726 50614
rect 154490 50058 154726 50294
rect 159610 54098 159846 54334
rect 159610 53778 159846 54014
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221050 414098 221286 414334
rect 221050 413778 221286 414014
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 215930 374378 216166 374614
rect 215930 374058 216166 374294
rect 210810 370658 211046 370894
rect 210810 370338 211046 370574
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 205690 330938 205926 331174
rect 205690 330618 205926 330854
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 200570 291218 200806 291454
rect 200570 290898 200806 291134
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 195450 237818 195686 238054
rect 195450 237498 195686 237734
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 190330 198098 190566 198334
rect 190330 197778 190566 198014
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 185210 158378 185446 158614
rect 185210 158058 185446 158294
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 180090 118658 180326 118894
rect 180090 118338 180326 118574
rect 174970 114938 175206 115174
rect 174970 114618 175206 114854
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 169850 75218 170086 75454
rect 169850 74898 170086 75134
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 164730 57818 164966 58054
rect 164730 57498 164966 57734
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 134010 21818 134246 22054
rect 134010 21498 134246 21734
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 144250 6938 144486 7174
rect 144250 6618 144486 6854
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 149370 10658 149606 10894
rect 149370 10338 149606 10574
rect 154490 14378 154726 14614
rect 154490 14058 154726 14294
rect 159610 18098 159846 18334
rect 159610 17778 159846 18014
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221050 378098 221286 378334
rect 221050 377778 221286 378014
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 215930 338378 216166 338614
rect 215930 338058 216166 338294
rect 210810 334658 211046 334894
rect 210810 334338 211046 334574
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 205690 294938 205926 295174
rect 205690 294618 205926 294854
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 200570 255218 200806 255454
rect 200570 254898 200806 255134
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 195450 201818 195686 202054
rect 195450 201498 195686 201734
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 190330 162098 190566 162334
rect 190330 161778 190566 162014
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 185210 122378 185446 122614
rect 185210 122058 185446 122294
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 180090 82658 180326 82894
rect 180090 82338 180326 82574
rect 174970 78938 175206 79174
rect 174970 78618 175206 78854
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 169850 39218 170086 39454
rect 169850 38898 170086 39134
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 164730 21818 164966 22054
rect 164730 21498 164966 21734
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221050 342098 221286 342334
rect 221050 341778 221286 342014
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 215930 302378 216166 302614
rect 215930 302058 216166 302294
rect 210810 298658 211046 298894
rect 210810 298338 211046 298574
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 205690 258938 205926 259174
rect 205690 258618 205926 258854
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 200570 219218 200806 219454
rect 200570 218898 200806 219134
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 195450 165818 195686 166054
rect 195450 165498 195686 165734
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 190330 126098 190566 126334
rect 190330 125778 190566 126014
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 185210 86378 185446 86614
rect 185210 86058 185446 86294
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 180090 46658 180326 46894
rect 180090 46338 180326 46574
rect 174970 42938 175206 43174
rect 174970 42618 175206 42854
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221050 306098 221286 306334
rect 221050 305778 221286 306014
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 215930 266378 216166 266614
rect 215930 266058 216166 266294
rect 210810 262658 211046 262894
rect 210810 262338 211046 262574
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 205690 222938 205926 223174
rect 205690 222618 205926 222854
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 200570 183218 200806 183454
rect 200570 182898 200806 183134
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 195450 129818 195686 130054
rect 195450 129498 195686 129734
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 190330 90098 190566 90334
rect 190330 89778 190566 90014
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 185210 50378 185446 50614
rect 185210 50058 185446 50294
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 180090 10658 180326 10894
rect 180090 10338 180326 10574
rect 174970 6938 175206 7174
rect 174970 6618 175206 6854
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221050 270098 221286 270334
rect 221050 269778 221286 270014
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 215930 230378 216166 230614
rect 215930 230058 216166 230294
rect 210810 226658 211046 226894
rect 210810 226338 211046 226574
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 205690 186938 205926 187174
rect 205690 186618 205926 186854
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 200570 147218 200806 147454
rect 200570 146898 200806 147134
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 195450 93818 195686 94054
rect 195450 93498 195686 93734
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 190330 54098 190566 54334
rect 190330 53778 190566 54014
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 185210 14378 185446 14614
rect 185210 14058 185446 14294
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221050 234098 221286 234334
rect 221050 233778 221286 234014
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 215930 194378 216166 194614
rect 215930 194058 216166 194294
rect 210810 190658 211046 190894
rect 210810 190338 211046 190574
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 205690 150938 205926 151174
rect 205690 150618 205926 150854
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 200570 111218 200806 111454
rect 200570 110898 200806 111134
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 195450 57818 195686 58054
rect 195450 57498 195686 57734
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 190330 18098 190566 18334
rect 190330 17778 190566 18014
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221050 198098 221286 198334
rect 221050 197778 221286 198014
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 215930 158378 216166 158614
rect 215930 158058 216166 158294
rect 210810 154658 211046 154894
rect 210810 154338 211046 154574
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 205690 114938 205926 115174
rect 205690 114618 205926 114854
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 200570 75218 200806 75454
rect 200570 74898 200806 75134
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 195450 21818 195686 22054
rect 195450 21498 195686 21734
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221050 162098 221286 162334
rect 221050 161778 221286 162014
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 215930 122378 216166 122614
rect 215930 122058 216166 122294
rect 210810 118658 211046 118894
rect 210810 118338 211046 118574
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 205690 78938 205926 79174
rect 205690 78618 205926 78854
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 200570 39218 200806 39454
rect 200570 38898 200806 39134
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221050 126098 221286 126334
rect 221050 125778 221286 126014
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 215930 86378 216166 86614
rect 215930 86058 216166 86294
rect 210810 82658 211046 82894
rect 210810 82338 211046 82574
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 205690 42938 205926 43174
rect 205690 42618 205926 42854
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221050 90098 221286 90334
rect 221050 89778 221286 90014
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 215930 50378 216166 50614
rect 215930 50058 216166 50294
rect 210810 46658 211046 46894
rect 210810 46338 211046 46574
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 205690 6938 205926 7174
rect 205690 6618 205926 6854
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221050 54098 221286 54334
rect 221050 53778 221286 54014
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 215930 14378 216166 14614
rect 215930 14058 216166 14294
rect 210810 10658 211046 10894
rect 210810 10338 211046 10574
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221050 18098 221286 18334
rect 221050 17778 221286 18014
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 226170 597818 226406 598054
rect 226170 597498 226406 597734
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 226170 561818 226406 562054
rect 226170 561498 226406 561734
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 232706 594098 232942 594334
rect 233026 594098 233262 594334
rect 232706 593778 232942 594014
rect 233026 593778 233262 594014
rect 231290 579218 231526 579454
rect 231290 578898 231526 579134
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 226170 525818 226406 526054
rect 226170 525498 226406 525734
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 240146 601538 240382 601774
rect 240466 601538 240702 601774
rect 240146 601218 240382 601454
rect 240466 601218 240702 601454
rect 236410 582938 236646 583174
rect 236410 582618 236646 582854
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 231290 543218 231526 543454
rect 231290 542898 231526 543134
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 226170 489818 226406 490054
rect 226170 489498 226406 489734
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 243866 605258 244102 605494
rect 244186 605258 244422 605494
rect 243866 604938 244102 605174
rect 244186 604938 244422 605174
rect 241530 586658 241766 586894
rect 241530 586338 241766 586574
rect 240146 565538 240382 565774
rect 240466 565538 240702 565774
rect 240146 565218 240382 565454
rect 240466 565218 240702 565454
rect 236410 546938 236646 547174
rect 236410 546618 236646 546854
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 231290 507218 231526 507454
rect 231290 506898 231526 507134
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 226170 453818 226406 454054
rect 226170 453498 226406 453734
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 251770 594098 252006 594334
rect 251770 593778 252006 594014
rect 246650 590378 246886 590614
rect 246650 590058 246886 590294
rect 243866 569258 244102 569494
rect 244186 569258 244422 569494
rect 243866 568938 244102 569174
rect 244186 568938 244422 569174
rect 241530 550658 241766 550894
rect 241530 550338 241766 550574
rect 240146 529538 240382 529774
rect 240466 529538 240702 529774
rect 240146 529218 240382 529454
rect 240466 529218 240702 529454
rect 236410 510938 236646 511174
rect 236410 510618 236646 510854
rect 232706 486098 232942 486334
rect 233026 486098 233262 486334
rect 232706 485778 232942 486014
rect 233026 485778 233262 486014
rect 231290 471218 231526 471454
rect 231290 470898 231526 471134
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 226170 417818 226406 418054
rect 226170 417498 226406 417734
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 256890 597818 257126 598054
rect 256890 597498 257126 597734
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 251770 558098 252006 558334
rect 251770 557778 252006 558014
rect 246650 554378 246886 554614
rect 246650 554058 246886 554294
rect 243866 533258 244102 533494
rect 244186 533258 244422 533494
rect 243866 532938 244102 533174
rect 244186 532938 244422 533174
rect 241530 514658 241766 514894
rect 241530 514338 241766 514574
rect 240146 493538 240382 493774
rect 240466 493538 240702 493774
rect 240146 493218 240382 493454
rect 240466 493218 240702 493454
rect 236410 474938 236646 475174
rect 236410 474618 236646 474854
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 231290 435218 231526 435454
rect 231290 434898 231526 435134
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 226170 381818 226406 382054
rect 226170 381498 226406 381734
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 256890 561818 257126 562054
rect 256890 561498 257126 561734
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 251770 522098 252006 522334
rect 251770 521778 252006 522014
rect 246650 518378 246886 518614
rect 246650 518058 246886 518294
rect 243866 497258 244102 497494
rect 244186 497258 244422 497494
rect 243866 496938 244102 497174
rect 244186 496938 244422 497174
rect 241530 478658 241766 478894
rect 241530 478338 241766 478574
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 236410 438938 236646 439174
rect 236410 438618 236646 438854
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 231290 399218 231526 399454
rect 231290 398898 231526 399134
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 226170 345818 226406 346054
rect 226170 345498 226406 345734
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 262010 579218 262246 579454
rect 262010 578898 262246 579134
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 256890 525818 257126 526054
rect 256890 525498 257126 525734
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 251770 486098 252006 486334
rect 251770 485778 252006 486014
rect 246650 482378 246886 482614
rect 246650 482058 246886 482294
rect 243866 461258 244102 461494
rect 244186 461258 244422 461494
rect 243866 460938 244102 461174
rect 244186 460938 244422 461174
rect 241530 442658 241766 442894
rect 241530 442338 241766 442574
rect 240146 421538 240382 421774
rect 240466 421538 240702 421774
rect 240146 421218 240382 421454
rect 240466 421218 240702 421454
rect 236410 402938 236646 403174
rect 236410 402618 236646 402854
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 231290 363218 231526 363454
rect 231290 362898 231526 363134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 226170 309818 226406 310054
rect 226170 309498 226406 309734
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 268706 594098 268942 594334
rect 269026 594098 269262 594334
rect 268706 593778 268942 594014
rect 269026 593778 269262 594014
rect 267130 582938 267366 583174
rect 267130 582618 267366 582854
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 262010 543218 262246 543454
rect 262010 542898 262246 543134
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 256890 489818 257126 490054
rect 256890 489498 257126 489734
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 251770 450098 252006 450334
rect 251770 449778 252006 450014
rect 246650 446378 246886 446614
rect 246650 446058 246886 446294
rect 243866 425258 244102 425494
rect 244186 425258 244422 425494
rect 243866 424938 244102 425174
rect 244186 424938 244422 425174
rect 241530 406658 241766 406894
rect 241530 406338 241766 406574
rect 240146 385538 240382 385774
rect 240466 385538 240702 385774
rect 240146 385218 240382 385454
rect 240466 385218 240702 385454
rect 236410 366938 236646 367174
rect 236410 366618 236646 366854
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 231290 327218 231526 327454
rect 231290 326898 231526 327134
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 226170 273818 226406 274054
rect 226170 273498 226406 273734
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 276146 601538 276382 601774
rect 276466 601538 276702 601774
rect 276146 601218 276382 601454
rect 276466 601218 276702 601454
rect 272250 586658 272486 586894
rect 272250 586338 272486 586574
rect 268706 558098 268942 558334
rect 269026 558098 269262 558334
rect 268706 557778 268942 558014
rect 269026 557778 269262 558014
rect 267130 546938 267366 547174
rect 267130 546618 267366 546854
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 262010 507218 262246 507454
rect 262010 506898 262246 507134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 256890 453818 257126 454054
rect 256890 453498 257126 453734
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 251770 414098 252006 414334
rect 251770 413778 252006 414014
rect 246650 410378 246886 410614
rect 246650 410058 246886 410294
rect 243866 389258 244102 389494
rect 244186 389258 244422 389494
rect 243866 388938 244102 389174
rect 244186 388938 244422 389174
rect 241530 370658 241766 370894
rect 241530 370338 241766 370574
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 236410 330938 236646 331174
rect 236410 330618 236646 330854
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 231290 291218 231526 291454
rect 231290 290898 231526 291134
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 226170 237818 226406 238054
rect 226170 237498 226406 237734
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 279866 605258 280102 605494
rect 280186 605258 280422 605494
rect 279866 604938 280102 605174
rect 280186 604938 280422 605174
rect 277370 590378 277606 590614
rect 277370 590058 277606 590294
rect 276146 565538 276382 565774
rect 276466 565538 276702 565774
rect 276146 565218 276382 565454
rect 276466 565218 276702 565454
rect 272250 550658 272486 550894
rect 272250 550338 272486 550574
rect 268706 522098 268942 522334
rect 269026 522098 269262 522334
rect 268706 521778 268942 522014
rect 269026 521778 269262 522014
rect 267130 510938 267366 511174
rect 267130 510618 267366 510854
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 262010 471218 262246 471454
rect 262010 470898 262246 471134
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 256890 417818 257126 418054
rect 256890 417498 257126 417734
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 251770 378098 252006 378334
rect 251770 377778 252006 378014
rect 246650 374378 246886 374614
rect 246650 374058 246886 374294
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 241530 334658 241766 334894
rect 241530 334338 241766 334574
rect 240146 313538 240382 313774
rect 240466 313538 240702 313774
rect 240146 313218 240382 313454
rect 240466 313218 240702 313454
rect 236410 294938 236646 295174
rect 236410 294618 236646 294854
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 231290 255218 231526 255454
rect 231290 254898 231526 255134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 226170 201818 226406 202054
rect 226170 201498 226406 201734
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 287610 597818 287846 598054
rect 287610 597498 287846 597734
rect 282490 594098 282726 594334
rect 282490 593778 282726 594014
rect 279866 569258 280102 569494
rect 280186 569258 280422 569494
rect 279866 568938 280102 569174
rect 280186 568938 280422 569174
rect 277370 554378 277606 554614
rect 277370 554058 277606 554294
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 272250 514658 272486 514894
rect 272250 514338 272486 514574
rect 268706 486098 268942 486334
rect 269026 486098 269262 486334
rect 268706 485778 268942 486014
rect 269026 485778 269262 486014
rect 267130 474938 267366 475174
rect 267130 474618 267366 474854
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 262010 435218 262246 435454
rect 262010 434898 262246 435134
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 256890 381818 257126 382054
rect 256890 381498 257126 381734
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 251770 342098 252006 342334
rect 251770 341778 252006 342014
rect 246650 338378 246886 338614
rect 246650 338058 246886 338294
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 241530 298658 241766 298894
rect 241530 298338 241766 298574
rect 240146 277538 240382 277774
rect 240466 277538 240702 277774
rect 240146 277218 240382 277454
rect 240466 277218 240702 277454
rect 236410 258938 236646 259174
rect 236410 258618 236646 258854
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 231290 219218 231526 219454
rect 231290 218898 231526 219134
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 226170 165818 226406 166054
rect 226170 165498 226406 165734
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 287610 561818 287846 562054
rect 287610 561498 287846 561734
rect 282490 558098 282726 558334
rect 282490 557778 282726 558014
rect 279866 533258 280102 533494
rect 280186 533258 280422 533494
rect 279866 532938 280102 533174
rect 280186 532938 280422 533174
rect 277370 518378 277606 518614
rect 277370 518058 277606 518294
rect 276146 493538 276382 493774
rect 276466 493538 276702 493774
rect 276146 493218 276382 493454
rect 276466 493218 276702 493454
rect 272250 478658 272486 478894
rect 272250 478338 272486 478574
rect 268706 450098 268942 450334
rect 269026 450098 269262 450334
rect 268706 449778 268942 450014
rect 269026 449778 269262 450014
rect 267130 438938 267366 439174
rect 267130 438618 267366 438854
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 262010 399218 262246 399454
rect 262010 398898 262246 399134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 256890 345818 257126 346054
rect 256890 345498 257126 345734
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 251770 306098 252006 306334
rect 251770 305778 252006 306014
rect 246650 302378 246886 302614
rect 246650 302058 246886 302294
rect 243866 281258 244102 281494
rect 244186 281258 244422 281494
rect 243866 280938 244102 281174
rect 244186 280938 244422 281174
rect 241530 262658 241766 262894
rect 241530 262338 241766 262574
rect 240146 241538 240382 241774
rect 240466 241538 240702 241774
rect 240146 241218 240382 241454
rect 240466 241218 240702 241454
rect 236410 222938 236646 223174
rect 236410 222618 236646 222854
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 231290 183218 231526 183454
rect 231290 182898 231526 183134
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 226170 129818 226406 130054
rect 226170 129498 226406 129734
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 292730 579218 292966 579454
rect 292730 578898 292966 579134
rect 297850 582938 298086 583174
rect 297850 582618 298086 582854
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 304706 630098 304942 630334
rect 305026 630098 305262 630334
rect 304706 629778 304942 630014
rect 305026 629778 305262 630014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 304706 594098 304942 594334
rect 305026 594098 305262 594334
rect 304706 593778 304942 594014
rect 305026 593778 305262 594014
rect 302970 586658 303206 586894
rect 302970 586338 303206 586574
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 287610 525818 287846 526054
rect 287610 525498 287846 525734
rect 282490 522098 282726 522334
rect 282490 521778 282726 522014
rect 279866 497258 280102 497494
rect 280186 497258 280422 497494
rect 279866 496938 280102 497174
rect 280186 496938 280422 497174
rect 277370 482378 277606 482614
rect 277370 482058 277606 482294
rect 276146 457538 276382 457774
rect 276466 457538 276702 457774
rect 276146 457218 276382 457454
rect 276466 457218 276702 457454
rect 272250 442658 272486 442894
rect 272250 442338 272486 442574
rect 268706 414098 268942 414334
rect 269026 414098 269262 414334
rect 268706 413778 268942 414014
rect 269026 413778 269262 414014
rect 267130 402938 267366 403174
rect 267130 402618 267366 402854
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 262010 363218 262246 363454
rect 262010 362898 262246 363134
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 256890 309818 257126 310054
rect 256890 309498 257126 309734
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 251770 270098 252006 270334
rect 251770 269778 252006 270014
rect 246650 266378 246886 266614
rect 246650 266058 246886 266294
rect 243866 245258 244102 245494
rect 244186 245258 244422 245494
rect 243866 244938 244102 245174
rect 244186 244938 244422 245174
rect 241530 226658 241766 226894
rect 241530 226338 241766 226574
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 236410 186938 236646 187174
rect 236410 186618 236646 186854
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 231290 147218 231526 147454
rect 231290 146898 231526 147134
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 226170 93818 226406 94054
rect 226170 93498 226406 93734
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 292730 543218 292966 543454
rect 292730 542898 292966 543134
rect 297850 546938 298086 547174
rect 297850 546618 298086 546854
rect 312146 601538 312382 601774
rect 312466 601538 312702 601774
rect 312146 601218 312382 601454
rect 312466 601218 312702 601454
rect 308090 590378 308326 590614
rect 308090 590058 308326 590294
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 302970 550658 303206 550894
rect 302970 550338 303206 550574
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 287610 489818 287846 490054
rect 287610 489498 287846 489734
rect 282490 486098 282726 486334
rect 282490 485778 282726 486014
rect 279866 461258 280102 461494
rect 280186 461258 280422 461494
rect 279866 460938 280102 461174
rect 280186 460938 280422 461174
rect 277370 446378 277606 446614
rect 277370 446058 277606 446294
rect 276146 421538 276382 421774
rect 276466 421538 276702 421774
rect 276146 421218 276382 421454
rect 276466 421218 276702 421454
rect 272250 406658 272486 406894
rect 272250 406338 272486 406574
rect 268706 378098 268942 378334
rect 269026 378098 269262 378334
rect 268706 377778 268942 378014
rect 269026 377778 269262 378014
rect 267130 366938 267366 367174
rect 267130 366618 267366 366854
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 262010 327218 262246 327454
rect 262010 326898 262246 327134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 256890 273818 257126 274054
rect 256890 273498 257126 273734
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 251770 234098 252006 234334
rect 251770 233778 252006 234014
rect 246650 230378 246886 230614
rect 246650 230058 246886 230294
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 241530 190658 241766 190894
rect 241530 190338 241766 190574
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 236410 150938 236646 151174
rect 236410 150618 236646 150854
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 231290 111218 231526 111454
rect 231290 110898 231526 111134
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 226170 57818 226406 58054
rect 226170 57498 226406 57734
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 292730 507218 292966 507454
rect 292730 506898 292966 507134
rect 297850 510938 298086 511174
rect 297850 510618 298086 510854
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 315866 605258 316102 605494
rect 316186 605258 316422 605494
rect 315866 604938 316102 605174
rect 316186 604938 316422 605174
rect 313210 594098 313446 594334
rect 313210 593778 313446 594014
rect 312146 565538 312382 565774
rect 312466 565538 312702 565774
rect 312146 565218 312382 565454
rect 312466 565218 312702 565454
rect 308090 554378 308326 554614
rect 308090 554058 308326 554294
rect 304706 522098 304942 522334
rect 305026 522098 305262 522334
rect 304706 521778 304942 522014
rect 305026 521778 305262 522014
rect 302970 514658 303206 514894
rect 302970 514338 303206 514574
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 287610 453818 287846 454054
rect 287610 453498 287846 453734
rect 282490 450098 282726 450334
rect 282490 449778 282726 450014
rect 279866 425258 280102 425494
rect 280186 425258 280422 425494
rect 279866 424938 280102 425174
rect 280186 424938 280422 425174
rect 277370 410378 277606 410614
rect 277370 410058 277606 410294
rect 276146 385538 276382 385774
rect 276466 385538 276702 385774
rect 276146 385218 276382 385454
rect 276466 385218 276702 385454
rect 272250 370658 272486 370894
rect 272250 370338 272486 370574
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 267130 330938 267366 331174
rect 267130 330618 267366 330854
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 262010 291218 262246 291454
rect 262010 290898 262246 291134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 256890 237818 257126 238054
rect 256890 237498 257126 237734
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 251770 198098 252006 198334
rect 251770 197778 252006 198014
rect 246650 194378 246886 194614
rect 246650 194058 246886 194294
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 241530 154658 241766 154894
rect 241530 154338 241766 154574
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 236410 114938 236646 115174
rect 236410 114618 236646 114854
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 231290 75218 231526 75454
rect 231290 74898 231526 75134
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 226170 21818 226406 22054
rect 226170 21498 226406 21734
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 292730 471218 292966 471454
rect 292730 470898 292966 471134
rect 297850 474938 298086 475174
rect 297850 474618 298086 474854
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 318330 597818 318566 598054
rect 318330 597498 318566 597734
rect 323450 579218 323686 579454
rect 323450 578898 323686 579134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 340706 630098 340942 630334
rect 341026 630098 341262 630334
rect 340706 629778 340942 630014
rect 341026 629778 341262 630014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 340706 594098 340942 594334
rect 341026 594098 341262 594334
rect 340706 593778 340942 594014
rect 341026 593778 341262 594014
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 333690 586658 333926 586894
rect 333690 586338 333926 586574
rect 338810 590378 339046 590614
rect 338810 590058 339046 590294
rect 343930 594098 344166 594334
rect 343930 593778 344166 594014
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 349050 597818 349286 598054
rect 349050 597498 349286 597734
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 364410 586658 364646 586894
rect 364410 586338 364646 586574
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 369530 590378 369766 590614
rect 369530 590058 369766 590294
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 374650 594098 374886 594334
rect 374650 593778 374886 594014
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 379770 597818 380006 598054
rect 379770 597498 380006 597734
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 395130 586658 395366 586894
rect 395130 586338 395366 586574
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 400250 590378 400486 590614
rect 400250 590058 400486 590294
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 405370 594098 405606 594334
rect 405370 593778 405606 594014
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 410490 597818 410726 598054
rect 410490 597498 410726 597734
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 328570 582938 328806 583174
rect 328570 582618 328806 582854
rect 359290 582938 359526 583174
rect 359290 582618 359526 582854
rect 390010 582938 390246 583174
rect 390010 582618 390246 582854
rect 420730 582938 420966 583174
rect 420730 582618 420966 582854
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 315866 569258 316102 569494
rect 316186 569258 316422 569494
rect 315866 568938 316102 569174
rect 316186 568938 316422 569174
rect 313210 558098 313446 558334
rect 313210 557778 313446 558014
rect 312146 529538 312382 529774
rect 312466 529538 312702 529774
rect 312146 529218 312382 529454
rect 312466 529218 312702 529454
rect 308090 518378 308326 518614
rect 308090 518058 308326 518294
rect 304706 486098 304942 486334
rect 305026 486098 305262 486334
rect 304706 485778 304942 486014
rect 305026 485778 305262 486014
rect 302970 478658 303206 478894
rect 302970 478338 303206 478574
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 287610 417818 287846 418054
rect 287610 417498 287846 417734
rect 282490 414098 282726 414334
rect 282490 413778 282726 414014
rect 279866 389258 280102 389494
rect 280186 389258 280422 389494
rect 279866 388938 280102 389174
rect 280186 388938 280422 389174
rect 277370 374378 277606 374614
rect 277370 374058 277606 374294
rect 276146 349538 276382 349774
rect 276466 349538 276702 349774
rect 276146 349218 276382 349454
rect 276466 349218 276702 349454
rect 272250 334658 272486 334894
rect 272250 334338 272486 334574
rect 268706 306098 268942 306334
rect 269026 306098 269262 306334
rect 268706 305778 268942 306014
rect 269026 305778 269262 306014
rect 267130 294938 267366 295174
rect 267130 294618 267366 294854
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 262010 255218 262246 255454
rect 262010 254898 262246 255134
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 256890 201818 257126 202054
rect 256890 201498 257126 201734
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 251770 162098 252006 162334
rect 251770 161778 252006 162014
rect 246650 158378 246886 158614
rect 246650 158058 246886 158294
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 241530 118658 241766 118894
rect 241530 118338 241766 118574
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 236410 78938 236646 79174
rect 236410 78618 236646 78854
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 231290 39218 231526 39454
rect 231290 38898 231526 39134
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 292730 435218 292966 435454
rect 292730 434898 292966 435134
rect 297850 438938 298086 439174
rect 297850 438618 298086 438854
rect 318330 561818 318566 562054
rect 318330 561498 318566 561734
rect 323450 543218 323686 543454
rect 323450 542898 323686 543134
rect 354170 579218 354406 579454
rect 354170 578898 354406 579134
rect 384890 579218 385126 579454
rect 384890 578898 385126 579134
rect 415610 579218 415846 579454
rect 415610 578898 415846 579134
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 430970 590378 431206 590614
rect 430970 590058 431206 590294
rect 425850 586658 426086 586894
rect 425850 586338 426086 586574
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 349050 561818 349286 562054
rect 349050 561498 349286 561734
rect 379770 561818 380006 562054
rect 379770 561498 380006 561734
rect 410490 561818 410726 562054
rect 410490 561498 410726 561734
rect 343930 558098 344166 558334
rect 343930 557778 344166 558014
rect 374650 558098 374886 558334
rect 374650 557778 374886 558014
rect 405370 558098 405606 558334
rect 405370 557778 405606 558014
rect 338810 554378 339046 554614
rect 338810 554058 339046 554294
rect 369530 554378 369766 554614
rect 369530 554058 369766 554294
rect 400250 554378 400486 554614
rect 400250 554058 400486 554294
rect 333690 550658 333926 550894
rect 333690 550338 333926 550574
rect 364410 550658 364646 550894
rect 364410 550338 364646 550574
rect 395130 550658 395366 550894
rect 395130 550338 395366 550574
rect 328570 546938 328806 547174
rect 328570 546618 328806 546854
rect 359290 546938 359526 547174
rect 359290 546618 359526 546854
rect 390010 546938 390246 547174
rect 390010 546618 390246 546854
rect 420730 546938 420966 547174
rect 420730 546618 420966 546854
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 315866 533258 316102 533494
rect 316186 533258 316422 533494
rect 315866 532938 316102 533174
rect 316186 532938 316422 533174
rect 313210 522098 313446 522334
rect 313210 521778 313446 522014
rect 312146 493538 312382 493774
rect 312466 493538 312702 493774
rect 312146 493218 312382 493454
rect 312466 493218 312702 493454
rect 308090 482378 308326 482614
rect 308090 482058 308326 482294
rect 304706 450098 304942 450334
rect 305026 450098 305262 450334
rect 304706 449778 304942 450014
rect 305026 449778 305262 450014
rect 302970 442658 303206 442894
rect 302970 442338 303206 442574
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 287610 381818 287846 382054
rect 287610 381498 287846 381734
rect 282490 378098 282726 378334
rect 282490 377778 282726 378014
rect 279866 353258 280102 353494
rect 280186 353258 280422 353494
rect 279866 352938 280102 353174
rect 280186 352938 280422 353174
rect 277370 338378 277606 338614
rect 277370 338058 277606 338294
rect 276146 313538 276382 313774
rect 276466 313538 276702 313774
rect 276146 313218 276382 313454
rect 276466 313218 276702 313454
rect 272250 298658 272486 298894
rect 272250 298338 272486 298574
rect 268706 270098 268942 270334
rect 269026 270098 269262 270334
rect 268706 269778 268942 270014
rect 269026 269778 269262 270014
rect 267130 258938 267366 259174
rect 267130 258618 267366 258854
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 262010 219218 262246 219454
rect 262010 218898 262246 219134
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 256890 165818 257126 166054
rect 256890 165498 257126 165734
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 251770 126098 252006 126334
rect 251770 125778 252006 126014
rect 246650 122378 246886 122614
rect 246650 122058 246886 122294
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 241530 82658 241766 82894
rect 241530 82338 241766 82574
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 236410 42938 236646 43174
rect 236410 42618 236646 42854
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 292730 399218 292966 399454
rect 292730 398898 292966 399134
rect 297850 402938 298086 403174
rect 297850 402618 298086 402854
rect 318330 525818 318566 526054
rect 318330 525498 318566 525734
rect 323450 507218 323686 507454
rect 323450 506898 323686 507134
rect 354170 543218 354406 543454
rect 354170 542898 354406 543134
rect 384890 543218 385126 543454
rect 384890 542898 385126 543134
rect 415610 543218 415846 543454
rect 415610 542898 415846 543134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 436090 594098 436326 594334
rect 436090 593778 436326 594014
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 430970 554378 431206 554614
rect 430970 554058 431206 554294
rect 425850 550658 426086 550894
rect 425850 550338 426086 550574
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 349050 525818 349286 526054
rect 349050 525498 349286 525734
rect 379770 525818 380006 526054
rect 379770 525498 380006 525734
rect 410490 525818 410726 526054
rect 410490 525498 410726 525734
rect 343930 522098 344166 522334
rect 343930 521778 344166 522014
rect 374650 522098 374886 522334
rect 374650 521778 374886 522014
rect 405370 522098 405606 522334
rect 405370 521778 405606 522014
rect 338810 518378 339046 518614
rect 338810 518058 339046 518294
rect 369530 518378 369766 518614
rect 369530 518058 369766 518294
rect 400250 518378 400486 518614
rect 400250 518058 400486 518294
rect 333690 514658 333926 514894
rect 333690 514338 333926 514574
rect 364410 514658 364646 514894
rect 364410 514338 364646 514574
rect 395130 514658 395366 514894
rect 395130 514338 395366 514574
rect 328570 510938 328806 511174
rect 328570 510618 328806 510854
rect 359290 510938 359526 511174
rect 359290 510618 359526 510854
rect 390010 510938 390246 511174
rect 390010 510618 390246 510854
rect 420730 510938 420966 511174
rect 420730 510618 420966 510854
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 315866 497258 316102 497494
rect 316186 497258 316422 497494
rect 315866 496938 316102 497174
rect 316186 496938 316422 497174
rect 313210 486098 313446 486334
rect 313210 485778 313446 486014
rect 312146 457538 312382 457774
rect 312466 457538 312702 457774
rect 312146 457218 312382 457454
rect 312466 457218 312702 457454
rect 308090 446378 308326 446614
rect 308090 446058 308326 446294
rect 304706 414098 304942 414334
rect 305026 414098 305262 414334
rect 304706 413778 304942 414014
rect 305026 413778 305262 414014
rect 302970 406658 303206 406894
rect 302970 406338 303206 406574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 287610 345818 287846 346054
rect 287610 345498 287846 345734
rect 282490 342098 282726 342334
rect 282490 341778 282726 342014
rect 279866 317258 280102 317494
rect 280186 317258 280422 317494
rect 279866 316938 280102 317174
rect 280186 316938 280422 317174
rect 277370 302378 277606 302614
rect 277370 302058 277606 302294
rect 276146 277538 276382 277774
rect 276466 277538 276702 277774
rect 276146 277218 276382 277454
rect 276466 277218 276702 277454
rect 272250 262658 272486 262894
rect 272250 262338 272486 262574
rect 268706 234098 268942 234334
rect 269026 234098 269262 234334
rect 268706 233778 268942 234014
rect 269026 233778 269262 234014
rect 267130 222938 267366 223174
rect 267130 222618 267366 222854
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 262010 183218 262246 183454
rect 262010 182898 262246 183134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 256890 129818 257126 130054
rect 256890 129498 257126 129734
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 251770 90098 252006 90334
rect 251770 89778 252006 90014
rect 246650 86378 246886 86614
rect 246650 86058 246886 86294
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 241530 46658 241766 46894
rect 241530 46338 241766 46574
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 236410 6938 236646 7174
rect 236410 6618 236646 6854
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 292730 363218 292966 363454
rect 292730 362898 292966 363134
rect 297850 366938 298086 367174
rect 297850 366618 298086 366854
rect 318330 489818 318566 490054
rect 318330 489498 318566 489734
rect 323450 471218 323686 471454
rect 323450 470898 323686 471134
rect 354170 507218 354406 507454
rect 354170 506898 354406 507134
rect 384890 507218 385126 507454
rect 384890 506898 385126 507134
rect 415610 507218 415846 507454
rect 415610 506898 415846 507134
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 441210 597818 441446 598054
rect 441210 597498 441446 597734
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 436090 558098 436326 558334
rect 436090 557778 436326 558014
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 430970 518378 431206 518614
rect 430970 518058 431206 518294
rect 425850 514658 426086 514894
rect 425850 514338 426086 514574
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 349050 489818 349286 490054
rect 349050 489498 349286 489734
rect 379770 489818 380006 490054
rect 379770 489498 380006 489734
rect 410490 489818 410726 490054
rect 410490 489498 410726 489734
rect 343930 486098 344166 486334
rect 343930 485778 344166 486014
rect 374650 486098 374886 486334
rect 374650 485778 374886 486014
rect 405370 486098 405606 486334
rect 405370 485778 405606 486014
rect 338810 482378 339046 482614
rect 338810 482058 339046 482294
rect 369530 482378 369766 482614
rect 369530 482058 369766 482294
rect 400250 482378 400486 482614
rect 400250 482058 400486 482294
rect 333690 478658 333926 478894
rect 333690 478338 333926 478574
rect 364410 478658 364646 478894
rect 364410 478338 364646 478574
rect 395130 478658 395366 478894
rect 395130 478338 395366 478574
rect 328570 474938 328806 475174
rect 328570 474618 328806 474854
rect 359290 474938 359526 475174
rect 359290 474618 359526 474854
rect 390010 474938 390246 475174
rect 390010 474618 390246 474854
rect 420730 474938 420966 475174
rect 420730 474618 420966 474854
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 315866 461258 316102 461494
rect 316186 461258 316422 461494
rect 315866 460938 316102 461174
rect 316186 460938 316422 461174
rect 313210 450098 313446 450334
rect 313210 449778 313446 450014
rect 312146 421538 312382 421774
rect 312466 421538 312702 421774
rect 312146 421218 312382 421454
rect 312466 421218 312702 421454
rect 308090 410378 308326 410614
rect 308090 410058 308326 410294
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 302970 370658 303206 370894
rect 302970 370338 303206 370574
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 287610 309818 287846 310054
rect 287610 309498 287846 309734
rect 282490 306098 282726 306334
rect 282490 305778 282726 306014
rect 279866 281258 280102 281494
rect 280186 281258 280422 281494
rect 279866 280938 280102 281174
rect 280186 280938 280422 281174
rect 277370 266378 277606 266614
rect 277370 266058 277606 266294
rect 276146 241538 276382 241774
rect 276466 241538 276702 241774
rect 276146 241218 276382 241454
rect 276466 241218 276702 241454
rect 272250 226658 272486 226894
rect 272250 226338 272486 226574
rect 268706 198098 268942 198334
rect 269026 198098 269262 198334
rect 268706 197778 268942 198014
rect 269026 197778 269262 198014
rect 267130 186938 267366 187174
rect 267130 186618 267366 186854
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 262010 147218 262246 147454
rect 262010 146898 262246 147134
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 256890 93818 257126 94054
rect 256890 93498 257126 93734
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 251770 54098 252006 54334
rect 251770 53778 252006 54014
rect 246650 50378 246886 50614
rect 246650 50058 246886 50294
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 241530 10658 241766 10894
rect 241530 10338 241766 10574
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 292730 327218 292966 327454
rect 292730 326898 292966 327134
rect 297850 330938 298086 331174
rect 297850 330618 298086 330854
rect 318330 453818 318566 454054
rect 318330 453498 318566 453734
rect 323450 435218 323686 435454
rect 323450 434898 323686 435134
rect 354170 471218 354406 471454
rect 354170 470898 354406 471134
rect 384890 471218 385126 471454
rect 384890 470898 385126 471134
rect 415610 471218 415846 471454
rect 415610 470898 415846 471134
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 441210 561818 441446 562054
rect 441210 561498 441446 561734
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 436090 522098 436326 522334
rect 436090 521778 436326 522014
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 430970 482378 431206 482614
rect 430970 482058 431206 482294
rect 425850 478658 426086 478894
rect 425850 478338 426086 478574
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 349050 453818 349286 454054
rect 349050 453498 349286 453734
rect 379770 453818 380006 454054
rect 379770 453498 380006 453734
rect 410490 453818 410726 454054
rect 410490 453498 410726 453734
rect 343930 450098 344166 450334
rect 343930 449778 344166 450014
rect 374650 450098 374886 450334
rect 374650 449778 374886 450014
rect 405370 450098 405606 450334
rect 405370 449778 405606 450014
rect 338810 446378 339046 446614
rect 338810 446058 339046 446294
rect 369530 446378 369766 446614
rect 369530 446058 369766 446294
rect 400250 446378 400486 446614
rect 400250 446058 400486 446294
rect 333690 442658 333926 442894
rect 333690 442338 333926 442574
rect 364410 442658 364646 442894
rect 364410 442338 364646 442574
rect 395130 442658 395366 442894
rect 395130 442338 395366 442574
rect 328570 438938 328806 439174
rect 328570 438618 328806 438854
rect 359290 438938 359526 439174
rect 359290 438618 359526 438854
rect 390010 438938 390246 439174
rect 390010 438618 390246 438854
rect 420730 438938 420966 439174
rect 420730 438618 420966 438854
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 315866 425258 316102 425494
rect 316186 425258 316422 425494
rect 315866 424938 316102 425174
rect 316186 424938 316422 425174
rect 313210 414098 313446 414334
rect 313210 413778 313446 414014
rect 312146 385538 312382 385774
rect 312466 385538 312702 385774
rect 312146 385218 312382 385454
rect 312466 385218 312702 385454
rect 308090 374378 308326 374614
rect 308090 374058 308326 374294
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 302970 334658 303206 334894
rect 302970 334338 303206 334574
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 287610 273818 287846 274054
rect 287610 273498 287846 273734
rect 282490 270098 282726 270334
rect 282490 269778 282726 270014
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 277370 230378 277606 230614
rect 277370 230058 277606 230294
rect 276146 205538 276382 205774
rect 276466 205538 276702 205774
rect 276146 205218 276382 205454
rect 276466 205218 276702 205454
rect 272250 190658 272486 190894
rect 272250 190338 272486 190574
rect 268706 162098 268942 162334
rect 269026 162098 269262 162334
rect 268706 161778 268942 162014
rect 269026 161778 269262 162014
rect 267130 150938 267366 151174
rect 267130 150618 267366 150854
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 262010 111218 262246 111454
rect 262010 110898 262246 111134
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 256890 57818 257126 58054
rect 256890 57498 257126 57734
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 251770 18098 252006 18334
rect 251770 17778 252006 18014
rect 246650 14378 246886 14614
rect 246650 14058 246886 14294
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 292730 291218 292966 291454
rect 292730 290898 292966 291134
rect 297850 294938 298086 295174
rect 297850 294618 298086 294854
rect 318330 417818 318566 418054
rect 318330 417498 318566 417734
rect 323450 399218 323686 399454
rect 323450 398898 323686 399134
rect 354170 435218 354406 435454
rect 354170 434898 354406 435134
rect 384890 435218 385126 435454
rect 384890 434898 385126 435134
rect 415610 435218 415846 435454
rect 415610 434898 415846 435134
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 446330 579218 446566 579454
rect 446330 578898 446566 579134
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 441210 525818 441446 526054
rect 441210 525498 441446 525734
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 436090 486098 436326 486334
rect 436090 485778 436326 486014
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 430970 446378 431206 446614
rect 430970 446058 431206 446294
rect 425850 442658 426086 442894
rect 425850 442338 426086 442574
rect 423866 425258 424102 425494
rect 424186 425258 424422 425494
rect 423866 424938 424102 425174
rect 424186 424938 424422 425174
rect 349050 417818 349286 418054
rect 349050 417498 349286 417734
rect 379770 417818 380006 418054
rect 379770 417498 380006 417734
rect 410490 417818 410726 418054
rect 410490 417498 410726 417734
rect 343930 414098 344166 414334
rect 343930 413778 344166 414014
rect 374650 414098 374886 414334
rect 374650 413778 374886 414014
rect 405370 414098 405606 414334
rect 405370 413778 405606 414014
rect 338810 410378 339046 410614
rect 338810 410058 339046 410294
rect 369530 410378 369766 410614
rect 369530 410058 369766 410294
rect 400250 410378 400486 410614
rect 400250 410058 400486 410294
rect 333690 406658 333926 406894
rect 333690 406338 333926 406574
rect 364410 406658 364646 406894
rect 364410 406338 364646 406574
rect 395130 406658 395366 406894
rect 395130 406338 395366 406574
rect 328570 402938 328806 403174
rect 328570 402618 328806 402854
rect 359290 402938 359526 403174
rect 359290 402618 359526 402854
rect 390010 402938 390246 403174
rect 390010 402618 390246 402854
rect 420730 402938 420966 403174
rect 420730 402618 420966 402854
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 315866 389258 316102 389494
rect 316186 389258 316422 389494
rect 315866 388938 316102 389174
rect 316186 388938 316422 389174
rect 313210 378098 313446 378334
rect 313210 377778 313446 378014
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 308090 338378 308326 338614
rect 308090 338058 308326 338294
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 302970 298658 303206 298894
rect 302970 298338 303206 298574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 287610 237818 287846 238054
rect 287610 237498 287846 237734
rect 282490 234098 282726 234334
rect 282490 233778 282726 234014
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 277370 194378 277606 194614
rect 277370 194058 277606 194294
rect 276146 169538 276382 169774
rect 276466 169538 276702 169774
rect 276146 169218 276382 169454
rect 276466 169218 276702 169454
rect 272250 154658 272486 154894
rect 272250 154338 272486 154574
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 267130 114938 267366 115174
rect 267130 114618 267366 114854
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 262010 75218 262246 75454
rect 262010 74898 262246 75134
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 256890 21818 257126 22054
rect 256890 21498 257126 21734
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 292730 255218 292966 255454
rect 292730 254898 292966 255134
rect 297850 258938 298086 259174
rect 297850 258618 298086 258854
rect 318330 381818 318566 382054
rect 318330 381498 318566 381734
rect 323450 363218 323686 363454
rect 323450 362898 323686 363134
rect 354170 399218 354406 399454
rect 354170 398898 354406 399134
rect 384890 399218 385126 399454
rect 384890 398898 385126 399134
rect 415610 399218 415846 399454
rect 415610 398898 415846 399134
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 451450 582938 451686 583174
rect 451450 582618 451686 582854
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 446330 543218 446566 543454
rect 446330 542898 446566 543134
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 441210 489818 441446 490054
rect 441210 489498 441446 489734
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 436090 450098 436326 450334
rect 436090 449778 436326 450014
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 430970 410378 431206 410614
rect 430970 410058 431206 410294
rect 425850 406658 426086 406894
rect 425850 406338 426086 406574
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 349050 381818 349286 382054
rect 349050 381498 349286 381734
rect 379770 381818 380006 382054
rect 379770 381498 380006 381734
rect 410490 381818 410726 382054
rect 410490 381498 410726 381734
rect 343930 378098 344166 378334
rect 343930 377778 344166 378014
rect 374650 378098 374886 378334
rect 374650 377778 374886 378014
rect 405370 378098 405606 378334
rect 405370 377778 405606 378014
rect 338810 374378 339046 374614
rect 338810 374058 339046 374294
rect 369530 374378 369766 374614
rect 369530 374058 369766 374294
rect 400250 374378 400486 374614
rect 400250 374058 400486 374294
rect 333690 370658 333926 370894
rect 333690 370338 333926 370574
rect 364410 370658 364646 370894
rect 364410 370338 364646 370574
rect 395130 370658 395366 370894
rect 395130 370338 395366 370574
rect 328570 366938 328806 367174
rect 328570 366618 328806 366854
rect 359290 366938 359526 367174
rect 359290 366618 359526 366854
rect 390010 366938 390246 367174
rect 390010 366618 390246 366854
rect 420730 366938 420966 367174
rect 420730 366618 420966 366854
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 313210 342098 313446 342334
rect 313210 341778 313446 342014
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 308090 302378 308326 302614
rect 308090 302058 308326 302294
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 302970 262658 303206 262894
rect 302970 262338 303206 262574
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 287610 201818 287846 202054
rect 287610 201498 287846 201734
rect 282490 198098 282726 198334
rect 282490 197778 282726 198014
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 277370 158378 277606 158614
rect 277370 158058 277606 158294
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 272250 118658 272486 118894
rect 272250 118338 272486 118574
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 267130 78938 267366 79174
rect 267130 78618 267366 78854
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 262010 39218 262246 39454
rect 262010 38898 262246 39134
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 292730 219218 292966 219454
rect 292730 218898 292966 219134
rect 297850 222938 298086 223174
rect 297850 222618 298086 222854
rect 318330 345818 318566 346054
rect 318330 345498 318566 345734
rect 323450 327218 323686 327454
rect 323450 326898 323686 327134
rect 354170 363218 354406 363454
rect 354170 362898 354406 363134
rect 384890 363218 385126 363454
rect 384890 362898 385126 363134
rect 415610 363218 415846 363454
rect 415610 362898 415846 363134
rect 456570 586658 456806 586894
rect 456570 586338 456806 586574
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 451450 546938 451686 547174
rect 451450 546618 451686 546854
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 446330 507218 446566 507454
rect 446330 506898 446566 507134
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 441210 453818 441446 454054
rect 441210 453498 441446 453734
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 436090 414098 436326 414334
rect 436090 413778 436326 414014
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 430970 374378 431206 374614
rect 430970 374058 431206 374294
rect 425850 370658 426086 370894
rect 425850 370338 426086 370574
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 349050 345818 349286 346054
rect 349050 345498 349286 345734
rect 379770 345818 380006 346054
rect 379770 345498 380006 345734
rect 410490 345818 410726 346054
rect 410490 345498 410726 345734
rect 343930 342098 344166 342334
rect 343930 341778 344166 342014
rect 374650 342098 374886 342334
rect 374650 341778 374886 342014
rect 405370 342098 405606 342334
rect 405370 341778 405606 342014
rect 338810 338378 339046 338614
rect 338810 338058 339046 338294
rect 369530 338378 369766 338614
rect 369530 338058 369766 338294
rect 400250 338378 400486 338614
rect 400250 338058 400486 338294
rect 333690 334658 333926 334894
rect 333690 334338 333926 334574
rect 364410 334658 364646 334894
rect 364410 334338 364646 334574
rect 395130 334658 395366 334894
rect 395130 334338 395366 334574
rect 328570 330938 328806 331174
rect 328570 330618 328806 330854
rect 359290 330938 359526 331174
rect 359290 330618 359526 330854
rect 390010 330938 390246 331174
rect 390010 330618 390246 330854
rect 420730 330938 420966 331174
rect 420730 330618 420966 330854
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 313210 306098 313446 306334
rect 313210 305778 313446 306014
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 308090 266378 308326 266614
rect 308090 266058 308326 266294
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 302970 226658 303206 226894
rect 302970 226338 303206 226574
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 287610 165818 287846 166054
rect 287610 165498 287846 165734
rect 282490 162098 282726 162334
rect 282490 161778 282726 162014
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 277370 122378 277606 122614
rect 277370 122058 277606 122294
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 272250 82658 272486 82894
rect 272250 82338 272486 82574
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 267130 42938 267366 43174
rect 267130 42618 267366 42854
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 292730 183218 292966 183454
rect 292730 182898 292966 183134
rect 297850 186938 298086 187174
rect 297850 186618 298086 186854
rect 318330 309818 318566 310054
rect 318330 309498 318566 309734
rect 323450 291218 323686 291454
rect 323450 290898 323686 291134
rect 354170 327218 354406 327454
rect 354170 326898 354406 327134
rect 384890 327218 385126 327454
rect 384890 326898 385126 327134
rect 415610 327218 415846 327454
rect 415610 326898 415846 327134
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 466810 594098 467046 594334
rect 466810 593778 467046 594014
rect 461690 590378 461926 590614
rect 461690 590058 461926 590294
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 456570 550658 456806 550894
rect 456570 550338 456806 550574
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 451450 510938 451686 511174
rect 451450 510618 451686 510854
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 446330 471218 446566 471454
rect 446330 470898 446566 471134
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 441210 417818 441446 418054
rect 441210 417498 441446 417734
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 436090 378098 436326 378334
rect 436090 377778 436326 378014
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 430970 338378 431206 338614
rect 430970 338058 431206 338294
rect 425850 334658 426086 334894
rect 425850 334338 426086 334574
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 349050 309818 349286 310054
rect 349050 309498 349286 309734
rect 379770 309818 380006 310054
rect 379770 309498 380006 309734
rect 410490 309818 410726 310054
rect 410490 309498 410726 309734
rect 343930 306098 344166 306334
rect 343930 305778 344166 306014
rect 374650 306098 374886 306334
rect 374650 305778 374886 306014
rect 405370 306098 405606 306334
rect 405370 305778 405606 306014
rect 338810 302378 339046 302614
rect 338810 302058 339046 302294
rect 369530 302378 369766 302614
rect 369530 302058 369766 302294
rect 400250 302378 400486 302614
rect 400250 302058 400486 302294
rect 333690 298658 333926 298894
rect 333690 298338 333926 298574
rect 364410 298658 364646 298894
rect 364410 298338 364646 298574
rect 395130 298658 395366 298894
rect 395130 298338 395366 298574
rect 328570 294938 328806 295174
rect 328570 294618 328806 294854
rect 359290 294938 359526 295174
rect 359290 294618 359526 294854
rect 390010 294938 390246 295174
rect 390010 294618 390246 294854
rect 420730 294938 420966 295174
rect 420730 294618 420966 294854
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 313210 270098 313446 270334
rect 313210 269778 313446 270014
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 308090 230378 308326 230614
rect 308090 230058 308326 230294
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 302970 190658 303206 190894
rect 302970 190338 303206 190574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 287610 129818 287846 130054
rect 287610 129498 287846 129734
rect 282490 126098 282726 126334
rect 282490 125778 282726 126014
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 277370 86378 277606 86614
rect 277370 86058 277606 86294
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 272250 46658 272486 46894
rect 272250 46338 272486 46574
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 267130 6938 267366 7174
rect 267130 6618 267366 6854
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 292730 147218 292966 147454
rect 292730 146898 292966 147134
rect 297850 150938 298086 151174
rect 297850 150618 298086 150854
rect 318330 273818 318566 274054
rect 318330 273498 318566 273734
rect 323450 255218 323686 255454
rect 323450 254898 323686 255134
rect 354170 291218 354406 291454
rect 354170 290898 354406 291134
rect 384890 291218 385126 291454
rect 384890 290898 385126 291134
rect 415610 291218 415846 291454
rect 415610 290898 415846 291134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 471930 597818 472166 598054
rect 471930 597498 472166 597734
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 466810 558098 467046 558334
rect 466810 557778 467046 558014
rect 461690 554378 461926 554614
rect 461690 554058 461926 554294
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 456570 514658 456806 514894
rect 456570 514338 456806 514574
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 451450 474938 451686 475174
rect 451450 474618 451686 474854
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 446330 435218 446566 435454
rect 446330 434898 446566 435134
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 441210 381818 441446 382054
rect 441210 381498 441446 381734
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 436090 342098 436326 342334
rect 436090 341778 436326 342014
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 430970 302378 431206 302614
rect 430970 302058 431206 302294
rect 425850 298658 426086 298894
rect 425850 298338 426086 298574
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 349050 273818 349286 274054
rect 349050 273498 349286 273734
rect 379770 273818 380006 274054
rect 379770 273498 380006 273734
rect 410490 273818 410726 274054
rect 410490 273498 410726 273734
rect 343930 270098 344166 270334
rect 343930 269778 344166 270014
rect 374650 270098 374886 270334
rect 374650 269778 374886 270014
rect 405370 270098 405606 270334
rect 405370 269778 405606 270014
rect 338810 266378 339046 266614
rect 338810 266058 339046 266294
rect 369530 266378 369766 266614
rect 369530 266058 369766 266294
rect 400250 266378 400486 266614
rect 400250 266058 400486 266294
rect 333690 262658 333926 262894
rect 333690 262338 333926 262574
rect 364410 262658 364646 262894
rect 364410 262338 364646 262574
rect 395130 262658 395366 262894
rect 395130 262338 395366 262574
rect 328570 258938 328806 259174
rect 328570 258618 328806 258854
rect 359290 258938 359526 259174
rect 359290 258618 359526 258854
rect 390010 258938 390246 259174
rect 390010 258618 390246 258854
rect 420730 258938 420966 259174
rect 420730 258618 420966 258854
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 313210 234098 313446 234334
rect 313210 233778 313446 234014
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 308090 194378 308326 194614
rect 308090 194058 308326 194294
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 302970 154658 303206 154894
rect 302970 154338 303206 154574
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 287610 93818 287846 94054
rect 287610 93498 287846 93734
rect 282490 90098 282726 90334
rect 282490 89778 282726 90014
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 277370 50378 277606 50614
rect 277370 50058 277606 50294
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 272250 10658 272486 10894
rect 272250 10338 272486 10574
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 292730 111218 292966 111454
rect 292730 110898 292966 111134
rect 297850 114938 298086 115174
rect 297850 114618 298086 114854
rect 318330 237818 318566 238054
rect 318330 237498 318566 237734
rect 323450 219218 323686 219454
rect 323450 218898 323686 219134
rect 354170 255218 354406 255454
rect 354170 254898 354406 255134
rect 384890 255218 385126 255454
rect 384890 254898 385126 255134
rect 415610 255218 415846 255454
rect 415610 254898 415846 255134
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 471930 561818 472166 562054
rect 471930 561498 472166 561734
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 466810 522098 467046 522334
rect 466810 521778 467046 522014
rect 461690 518378 461926 518614
rect 461690 518058 461926 518294
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 456570 478658 456806 478894
rect 456570 478338 456806 478574
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 451450 438938 451686 439174
rect 451450 438618 451686 438854
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 446330 399218 446566 399454
rect 446330 398898 446566 399134
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 441210 345818 441446 346054
rect 441210 345498 441446 345734
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 436090 306098 436326 306334
rect 436090 305778 436326 306014
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 430970 266378 431206 266614
rect 430970 266058 431206 266294
rect 425850 262658 426086 262894
rect 425850 262338 426086 262574
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 349050 237818 349286 238054
rect 349050 237498 349286 237734
rect 379770 237818 380006 238054
rect 379770 237498 380006 237734
rect 410490 237818 410726 238054
rect 410490 237498 410726 237734
rect 343930 234098 344166 234334
rect 343930 233778 344166 234014
rect 374650 234098 374886 234334
rect 374650 233778 374886 234014
rect 405370 234098 405606 234334
rect 405370 233778 405606 234014
rect 338810 230378 339046 230614
rect 338810 230058 339046 230294
rect 369530 230378 369766 230614
rect 369530 230058 369766 230294
rect 400250 230378 400486 230614
rect 400250 230058 400486 230294
rect 333690 226658 333926 226894
rect 333690 226338 333926 226574
rect 364410 226658 364646 226894
rect 364410 226338 364646 226574
rect 395130 226658 395366 226894
rect 395130 226338 395366 226574
rect 328570 222938 328806 223174
rect 328570 222618 328806 222854
rect 359290 222938 359526 223174
rect 359290 222618 359526 222854
rect 390010 222938 390246 223174
rect 390010 222618 390246 222854
rect 420730 222938 420966 223174
rect 420730 222618 420966 222854
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 313210 198098 313446 198334
rect 313210 197778 313446 198014
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 308090 158378 308326 158614
rect 308090 158058 308326 158294
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 302970 118658 303206 118894
rect 302970 118338 303206 118574
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 287610 57818 287846 58054
rect 287610 57498 287846 57734
rect 282490 54098 282726 54334
rect 282490 53778 282726 54014
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 277370 14378 277606 14614
rect 277370 14058 277606 14294
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 292730 75218 292966 75454
rect 292730 74898 292966 75134
rect 297850 78938 298086 79174
rect 297850 78618 298086 78854
rect 318330 201818 318566 202054
rect 318330 201498 318566 201734
rect 323450 183218 323686 183454
rect 323450 182898 323686 183134
rect 354170 219218 354406 219454
rect 354170 218898 354406 219134
rect 384890 219218 385126 219454
rect 384890 218898 385126 219134
rect 415610 219218 415846 219454
rect 415610 218898 415846 219134
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 477050 579218 477286 579454
rect 477050 578898 477286 579134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 471930 525818 472166 526054
rect 471930 525498 472166 525734
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 466810 486098 467046 486334
rect 466810 485778 467046 486014
rect 461690 482378 461926 482614
rect 461690 482058 461926 482294
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 456570 442658 456806 442894
rect 456570 442338 456806 442574
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 451450 402938 451686 403174
rect 451450 402618 451686 402854
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 446330 363218 446566 363454
rect 446330 362898 446566 363134
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441210 309818 441446 310054
rect 441210 309498 441446 309734
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 436090 270098 436326 270334
rect 436090 269778 436326 270014
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 430970 230378 431206 230614
rect 430970 230058 431206 230294
rect 425850 226658 426086 226894
rect 425850 226338 426086 226574
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 349050 201818 349286 202054
rect 349050 201498 349286 201734
rect 379770 201818 380006 202054
rect 379770 201498 380006 201734
rect 410490 201818 410726 202054
rect 410490 201498 410726 201734
rect 343930 198098 344166 198334
rect 343930 197778 344166 198014
rect 374650 198098 374886 198334
rect 374650 197778 374886 198014
rect 338810 194378 339046 194614
rect 338810 194058 339046 194294
rect 369530 194378 369766 194614
rect 369530 194058 369766 194294
rect 400250 194195 400486 194431
rect 333690 190658 333926 190894
rect 333690 190338 333926 190574
rect 364410 190658 364646 190894
rect 364410 190338 364646 190574
rect 395130 190658 395366 190894
rect 395130 190338 395366 190574
rect 328570 186938 328806 187174
rect 328570 186618 328806 186854
rect 359290 186938 359526 187174
rect 359290 186618 359526 186854
rect 390010 186938 390246 187174
rect 390010 186618 390246 186854
rect 420730 186938 420966 187174
rect 420730 186618 420966 186854
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 313210 162098 313446 162334
rect 313210 161778 313446 162014
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 308090 122378 308326 122614
rect 308090 122058 308326 122294
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 302970 82658 303206 82894
rect 302970 82338 303206 82574
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 287610 21818 287846 22054
rect 287610 21498 287846 21734
rect 282490 18098 282726 18334
rect 282490 17778 282726 18014
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 292730 39218 292966 39454
rect 292730 38898 292966 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 297850 42938 298086 43174
rect 297850 42618 298086 42854
rect 318330 165818 318566 166054
rect 318330 165498 318566 165734
rect 323450 147218 323686 147454
rect 323450 146898 323686 147134
rect 354170 183218 354406 183454
rect 354170 182898 354406 183134
rect 384890 183218 385126 183454
rect 384890 182898 385126 183134
rect 415610 183218 415846 183454
rect 415610 182898 415846 183134
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 482170 582938 482406 583174
rect 482170 582618 482406 582854
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 477050 543218 477286 543454
rect 477050 542898 477286 543134
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 471930 489818 472166 490054
rect 471930 489498 472166 489734
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 466810 450098 467046 450334
rect 466810 449778 467046 450014
rect 461690 446378 461926 446614
rect 461690 446058 461926 446294
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 456570 406658 456806 406894
rect 456570 406338 456806 406574
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 451450 366938 451686 367174
rect 451450 366618 451686 366854
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 446330 327218 446566 327454
rect 446330 326898 446566 327134
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 441210 273818 441446 274054
rect 441210 273498 441446 273734
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 436090 234098 436326 234334
rect 436090 233778 436326 234014
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 430970 194378 431206 194614
rect 430970 194058 431206 194294
rect 425850 190658 426086 190894
rect 425850 190338 426086 190574
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 349050 165818 349286 166054
rect 349050 165498 349286 165734
rect 379770 165818 380006 166054
rect 379770 165498 380006 165734
rect 410490 165818 410726 166054
rect 410490 165498 410726 165734
rect 343930 162098 344166 162334
rect 343930 161778 344166 162014
rect 374650 162098 374886 162334
rect 374650 161778 374886 162014
rect 405370 162098 405606 162334
rect 405370 161778 405606 162014
rect 338810 158378 339046 158614
rect 338810 158058 339046 158294
rect 369530 158378 369766 158614
rect 369530 158058 369766 158294
rect 400250 158378 400486 158614
rect 400250 158058 400486 158294
rect 333690 154658 333926 154894
rect 333690 154338 333926 154574
rect 364410 154658 364646 154894
rect 364410 154338 364646 154574
rect 395130 154658 395366 154894
rect 395130 154338 395366 154574
rect 328570 150938 328806 151174
rect 328570 150618 328806 150854
rect 359290 150938 359526 151174
rect 359290 150618 359526 150854
rect 390010 150938 390246 151174
rect 390010 150618 390246 150854
rect 420730 150938 420966 151174
rect 420730 150618 420966 150854
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 313210 126098 313446 126334
rect 313210 125778 313446 126014
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 308090 86378 308326 86614
rect 308090 86058 308326 86294
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 302970 46658 303206 46894
rect 302970 46338 303206 46574
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 297850 6938 298086 7174
rect 297850 6618 298086 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 318330 129818 318566 130054
rect 318330 129498 318566 129734
rect 323450 111218 323686 111454
rect 323450 110898 323686 111134
rect 354170 147218 354406 147454
rect 354170 146898 354406 147134
rect 384890 147218 385126 147454
rect 384890 146898 385126 147134
rect 415610 147218 415846 147454
rect 415610 146898 415846 147134
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 495866 641258 496102 641494
rect 496186 641258 496422 641494
rect 495866 640938 496102 641174
rect 496186 640938 496422 641174
rect 495866 605258 496102 605494
rect 496186 605258 496422 605494
rect 495866 604938 496102 605174
rect 496186 604938 496422 605174
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 487290 586658 487526 586894
rect 487290 586338 487526 586574
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 482170 546938 482406 547174
rect 482170 546618 482406 546854
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 477050 507218 477286 507454
rect 477050 506898 477286 507134
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 471930 453818 472166 454054
rect 471930 453498 472166 453734
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 466810 414098 467046 414334
rect 466810 413778 467046 414014
rect 461690 410378 461926 410614
rect 461690 410058 461926 410294
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 456570 370658 456806 370894
rect 456570 370338 456806 370574
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 451450 330938 451686 331174
rect 451450 330618 451686 330854
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 446330 291218 446566 291454
rect 446330 290898 446566 291134
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 441210 237818 441446 238054
rect 441210 237498 441446 237734
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 436090 198098 436326 198334
rect 436090 197778 436326 198014
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 430970 158378 431206 158614
rect 430970 158058 431206 158294
rect 425850 154658 426086 154894
rect 425850 154338 426086 154574
rect 423866 137258 424102 137494
rect 424186 137258 424422 137494
rect 423866 136938 424102 137174
rect 424186 136938 424422 137174
rect 349050 129818 349286 130054
rect 349050 129498 349286 129734
rect 379770 129818 380006 130054
rect 379770 129498 380006 129734
rect 410490 129818 410726 130054
rect 410490 129498 410726 129734
rect 343930 126098 344166 126334
rect 343930 125778 344166 126014
rect 374650 126098 374886 126334
rect 374650 125778 374886 126014
rect 405370 126098 405606 126334
rect 405370 125778 405606 126014
rect 338810 122378 339046 122614
rect 338810 122058 339046 122294
rect 369530 122378 369766 122614
rect 369530 122058 369766 122294
rect 400250 122378 400486 122614
rect 400250 122058 400486 122294
rect 333690 118658 333926 118894
rect 333690 118338 333926 118574
rect 364410 118658 364646 118894
rect 364410 118338 364646 118574
rect 395130 118658 395366 118894
rect 395130 118338 395366 118574
rect 328570 114938 328806 115174
rect 328570 114618 328806 114854
rect 359290 114938 359526 115174
rect 359290 114618 359526 114854
rect 390010 114938 390246 115174
rect 390010 114618 390246 114854
rect 420730 114938 420966 115174
rect 420730 114618 420966 114854
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 313210 90098 313446 90334
rect 313210 89778 313446 90014
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 308090 50378 308326 50614
rect 308090 50058 308326 50294
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 302970 10658 303206 10894
rect 302970 10338 303206 10574
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 318330 93818 318566 94054
rect 318330 93498 318566 93734
rect 323450 75218 323686 75454
rect 323450 74898 323686 75134
rect 354170 111218 354406 111454
rect 354170 110898 354406 111134
rect 384890 111218 385126 111454
rect 384890 110898 385126 111134
rect 415610 111218 415846 111454
rect 415610 110898 415846 111134
rect 492410 590378 492646 590614
rect 492410 590058 492646 590294
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 487290 550658 487526 550894
rect 487290 550338 487526 550574
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 482170 510938 482406 511174
rect 482170 510618 482406 510854
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 477050 471218 477286 471454
rect 477050 470898 477286 471134
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 471930 417818 472166 418054
rect 471930 417498 472166 417734
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 466810 378098 467046 378334
rect 466810 377778 467046 378014
rect 461690 374378 461926 374614
rect 461690 374058 461926 374294
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 456570 334658 456806 334894
rect 456570 334338 456806 334574
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 451450 294938 451686 295174
rect 451450 294618 451686 294854
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 446330 255218 446566 255454
rect 446330 254898 446566 255134
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 441210 201818 441446 202054
rect 441210 201498 441446 201734
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 436090 162098 436326 162334
rect 436090 161778 436326 162014
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 430970 122378 431206 122614
rect 430970 122058 431206 122294
rect 425850 118658 426086 118894
rect 425850 118338 426086 118574
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 349050 93818 349286 94054
rect 349050 93498 349286 93734
rect 379770 93818 380006 94054
rect 379770 93498 380006 93734
rect 410490 93818 410726 94054
rect 410490 93498 410726 93734
rect 343930 90098 344166 90334
rect 343930 89778 344166 90014
rect 374650 90098 374886 90334
rect 374650 89778 374886 90014
rect 405370 90098 405606 90334
rect 405370 89778 405606 90014
rect 338810 86378 339046 86614
rect 338810 86058 339046 86294
rect 369530 86378 369766 86614
rect 369530 86058 369766 86294
rect 400250 86378 400486 86614
rect 400250 86058 400486 86294
rect 333690 82658 333926 82894
rect 333690 82338 333926 82574
rect 364410 82658 364646 82894
rect 364410 82338 364646 82574
rect 395130 82658 395366 82894
rect 395130 82338 395366 82574
rect 328570 78938 328806 79174
rect 328570 78618 328806 78854
rect 359290 78938 359526 79174
rect 359290 78618 359526 78854
rect 390010 78938 390246 79174
rect 390010 78618 390246 78854
rect 420730 78938 420966 79174
rect 420730 78618 420966 78854
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 313210 54098 313446 54334
rect 313210 53778 313446 54014
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 308090 14378 308326 14614
rect 308090 14058 308326 14294
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 318330 57818 318566 58054
rect 318330 57498 318566 57734
rect 323450 39218 323686 39454
rect 323450 38898 323686 39134
rect 354170 75218 354406 75454
rect 354170 74898 354406 75134
rect 384890 75218 385126 75454
rect 384890 74898 385126 75134
rect 415610 75218 415846 75454
rect 415610 74898 415846 75134
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 502650 597818 502886 598054
rect 502650 597498 502886 597734
rect 497530 594098 497766 594334
rect 497530 593778 497766 594014
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 492410 554378 492646 554614
rect 492410 554058 492646 554294
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 487290 514658 487526 514894
rect 487290 514338 487526 514574
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 482170 474938 482406 475174
rect 482170 474618 482406 474854
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 477050 435218 477286 435454
rect 477050 434898 477286 435134
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 471930 381818 472166 382054
rect 471930 381498 472166 381734
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 466810 342098 467046 342334
rect 466810 341778 467046 342014
rect 461690 338378 461926 338614
rect 461690 338058 461926 338294
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 456570 298658 456806 298894
rect 456570 298338 456806 298574
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 451450 258938 451686 259174
rect 451450 258618 451686 258854
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 446330 219218 446566 219454
rect 446330 218898 446566 219134
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 441210 165818 441446 166054
rect 441210 165498 441446 165734
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 436090 126098 436326 126334
rect 436090 125778 436326 126014
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 430970 86378 431206 86614
rect 430970 86058 431206 86294
rect 425850 82658 426086 82894
rect 425850 82338 426086 82574
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 349050 57818 349286 58054
rect 349050 57498 349286 57734
rect 379770 57818 380006 58054
rect 379770 57498 380006 57734
rect 410490 57818 410726 58054
rect 410490 57498 410726 57734
rect 343930 54098 344166 54334
rect 343930 53778 344166 54014
rect 374650 54098 374886 54334
rect 374650 53778 374886 54014
rect 405370 54098 405606 54334
rect 405370 53778 405606 54014
rect 338810 50378 339046 50614
rect 338810 50058 339046 50294
rect 369530 50378 369766 50614
rect 369530 50058 369766 50294
rect 400250 50378 400486 50614
rect 400250 50058 400486 50294
rect 333690 46658 333926 46894
rect 333690 46338 333926 46574
rect 364410 46658 364646 46894
rect 364410 46338 364646 46574
rect 395130 46658 395366 46894
rect 395130 46338 395366 46574
rect 328570 42938 328806 43174
rect 328570 42618 328806 42854
rect 359290 42938 359526 43174
rect 359290 42618 359526 42854
rect 390010 42938 390246 43174
rect 390010 42618 390246 42854
rect 420730 42938 420966 43174
rect 420730 42618 420966 42854
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 313210 18098 313446 18334
rect 313210 17778 313446 18014
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 318330 21818 318566 22054
rect 318330 21498 318566 21734
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 354170 39218 354406 39454
rect 354170 38898 354406 39134
rect 384890 39218 385126 39454
rect 384890 38898 385126 39134
rect 415610 39218 415846 39454
rect 415610 38898 415846 39134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 502650 561818 502886 562054
rect 502650 561498 502886 561734
rect 497530 558098 497766 558334
rect 497530 557778 497766 558014
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 492410 518378 492646 518614
rect 492410 518058 492646 518294
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 487290 478658 487526 478894
rect 487290 478338 487526 478574
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 482170 438938 482406 439174
rect 482170 438618 482406 438854
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 477050 399218 477286 399454
rect 477050 398898 477286 399134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 471930 345818 472166 346054
rect 471930 345498 472166 345734
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 466810 306098 467046 306334
rect 466810 305778 467046 306014
rect 461690 302378 461926 302614
rect 461690 302058 461926 302294
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 456570 262658 456806 262894
rect 456570 262338 456806 262574
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 451450 222938 451686 223174
rect 451450 222618 451686 222854
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 446330 183218 446566 183454
rect 446330 182898 446566 183134
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 441210 129818 441446 130054
rect 441210 129498 441446 129734
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 436090 90098 436326 90334
rect 436090 89778 436326 90014
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 430970 50378 431206 50614
rect 430970 50058 431206 50294
rect 425850 46658 426086 46894
rect 425850 46338 426086 46574
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 349050 21818 349286 22054
rect 349050 21498 349286 21734
rect 379770 21818 380006 22054
rect 379770 21498 380006 21734
rect 410490 21818 410726 22054
rect 410490 21498 410726 21734
rect 343930 18098 344166 18334
rect 343930 17778 344166 18014
rect 374650 18098 374886 18334
rect 374650 17778 374886 18014
rect 405370 18098 405606 18334
rect 405370 17778 405606 18014
rect 338810 14378 339046 14614
rect 338810 14058 339046 14294
rect 369530 14378 369766 14614
rect 369530 14058 369766 14294
rect 400250 14378 400486 14614
rect 400250 14058 400486 14294
rect 333690 10658 333926 10894
rect 333690 10338 333926 10574
rect 364410 10658 364646 10894
rect 364410 10338 364646 10574
rect 395130 10658 395366 10894
rect 395130 10338 395366 10574
rect 328570 6938 328806 7174
rect 328570 6618 328806 6854
rect 359290 6938 359526 7174
rect 359290 6618 359526 6854
rect 390010 6938 390246 7174
rect 390010 6618 390246 6854
rect 420730 6938 420966 7174
rect 420730 6618 420966 6854
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 507770 579218 508006 579454
rect 507770 578898 508006 579134
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 502650 525818 502886 526054
rect 502650 525498 502886 525734
rect 497530 522098 497766 522334
rect 497530 521778 497766 522014
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 492410 482378 492646 482614
rect 492410 482058 492646 482294
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 487290 442658 487526 442894
rect 487290 442338 487526 442574
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 482170 402938 482406 403174
rect 482170 402618 482406 402854
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 477050 363218 477286 363454
rect 477050 362898 477286 363134
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 471930 309818 472166 310054
rect 471930 309498 472166 309734
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 466810 270098 467046 270334
rect 466810 269778 467046 270014
rect 461690 266378 461926 266614
rect 461690 266058 461926 266294
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 456570 226658 456806 226894
rect 456570 226338 456806 226574
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 451450 186938 451686 187174
rect 451450 186618 451686 186854
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 446330 147218 446566 147454
rect 446330 146898 446566 147134
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 441210 93818 441446 94054
rect 441210 93498 441446 93734
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 436090 54098 436326 54334
rect 436090 53778 436326 54014
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 430970 14378 431206 14614
rect 430970 14058 431206 14294
rect 425850 10658 426086 10894
rect 425850 10338 426086 10574
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 507770 543218 508006 543454
rect 507770 542898 508006 543134
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 502650 489818 502886 490054
rect 502650 489498 502886 489734
rect 497530 486098 497766 486334
rect 497530 485778 497766 486014
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 492410 446378 492646 446614
rect 492410 446058 492646 446294
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 487290 406658 487526 406894
rect 487290 406338 487526 406574
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 482170 366938 482406 367174
rect 482170 366618 482406 366854
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 477050 327218 477286 327454
rect 477050 326898 477286 327134
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 471930 273818 472166 274054
rect 471930 273498 472166 273734
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 466810 234098 467046 234334
rect 466810 233778 467046 234014
rect 461690 230378 461926 230614
rect 461690 230058 461926 230294
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 456570 190658 456806 190894
rect 456570 190338 456806 190574
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 451450 150938 451686 151174
rect 451450 150618 451686 150854
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 446330 111218 446566 111454
rect 446330 110898 446566 111134
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 441210 57818 441446 58054
rect 441210 57498 441446 57734
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 436090 18098 436326 18334
rect 436090 17778 436326 18014
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 507770 507218 508006 507454
rect 507770 506898 508006 507134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 502650 453818 502886 454054
rect 502650 453498 502886 453734
rect 497530 450098 497766 450334
rect 497530 449778 497766 450014
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 492410 410378 492646 410614
rect 492410 410058 492646 410294
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 487290 370658 487526 370894
rect 487290 370338 487526 370574
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 482170 330938 482406 331174
rect 482170 330618 482406 330854
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 477050 291218 477286 291454
rect 477050 290898 477286 291134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 471930 237818 472166 238054
rect 471930 237498 472166 237734
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 466810 198098 467046 198334
rect 466810 197778 467046 198014
rect 461690 194378 461926 194614
rect 461690 194058 461926 194294
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 456570 154658 456806 154894
rect 456570 154338 456806 154574
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 451450 114938 451686 115174
rect 451450 114618 451686 114854
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 446330 75218 446566 75454
rect 446330 74898 446566 75134
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 441210 21818 441446 22054
rect 441210 21498 441446 21734
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 507770 471218 508006 471454
rect 507770 470898 508006 471134
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 502650 417818 502886 418054
rect 502650 417498 502886 417734
rect 497530 414098 497766 414334
rect 497530 413778 497766 414014
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 492410 374378 492646 374614
rect 492410 374058 492646 374294
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 487290 334658 487526 334894
rect 487290 334338 487526 334574
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 482170 294938 482406 295174
rect 482170 294618 482406 294854
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 477050 255218 477286 255454
rect 477050 254898 477286 255134
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 471930 201818 472166 202054
rect 471930 201498 472166 201734
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 466810 162098 467046 162334
rect 466810 161778 467046 162014
rect 461690 158378 461926 158614
rect 461690 158058 461926 158294
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 456570 118658 456806 118894
rect 456570 118338 456806 118574
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 451450 78938 451686 79174
rect 451450 78618 451686 78854
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 446330 39218 446566 39454
rect 446330 38898 446566 39134
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 507770 435218 508006 435454
rect 507770 434898 508006 435134
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 502650 381818 502886 382054
rect 502650 381498 502886 381734
rect 497530 378098 497766 378334
rect 497530 377778 497766 378014
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 492410 338378 492646 338614
rect 492410 338058 492646 338294
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 487290 298658 487526 298894
rect 487290 298338 487526 298574
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 482170 258938 482406 259174
rect 482170 258618 482406 258854
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 477050 219218 477286 219454
rect 477050 218898 477286 219134
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 471930 165818 472166 166054
rect 471930 165498 472166 165734
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 466810 126098 467046 126334
rect 466810 125778 467046 126014
rect 461690 122378 461926 122614
rect 461690 122058 461926 122294
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 456570 82658 456806 82894
rect 456570 82338 456806 82574
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 451450 42938 451686 43174
rect 451450 42618 451686 42854
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 507770 399218 508006 399454
rect 507770 398898 508006 399134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 502650 345818 502886 346054
rect 502650 345498 502886 345734
rect 497530 342098 497766 342334
rect 497530 341778 497766 342014
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 492410 302378 492646 302614
rect 492410 302058 492646 302294
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 487290 262658 487526 262894
rect 487290 262338 487526 262574
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 482170 222938 482406 223174
rect 482170 222618 482406 222854
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 477050 183218 477286 183454
rect 477050 182898 477286 183134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 471930 129818 472166 130054
rect 471930 129498 472166 129734
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 466810 90098 467046 90334
rect 466810 89778 467046 90014
rect 461690 86378 461926 86614
rect 461690 86058 461926 86294
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 456570 46658 456806 46894
rect 456570 46338 456806 46574
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 451450 6938 451686 7174
rect 451450 6618 451686 6854
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 507770 363218 508006 363454
rect 507770 362898 508006 363134
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 502650 309818 502886 310054
rect 502650 309498 502886 309734
rect 497530 306098 497766 306334
rect 497530 305778 497766 306014
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 492410 266378 492646 266614
rect 492410 266058 492646 266294
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 487290 226658 487526 226894
rect 487290 226338 487526 226574
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 482170 186938 482406 187174
rect 482170 186618 482406 186854
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 477050 147218 477286 147454
rect 477050 146898 477286 147134
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 471930 93818 472166 94054
rect 471930 93498 472166 93734
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 466810 54098 467046 54334
rect 466810 53778 467046 54014
rect 461690 50378 461926 50614
rect 461690 50058 461926 50294
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 456570 10658 456806 10894
rect 456570 10338 456806 10574
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 507770 327218 508006 327454
rect 507770 326898 508006 327134
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 502650 273818 502886 274054
rect 502650 273498 502886 273734
rect 497530 270098 497766 270334
rect 497530 269778 497766 270014
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 492410 230378 492646 230614
rect 492410 230058 492646 230294
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 487290 190658 487526 190894
rect 487290 190338 487526 190574
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 482170 150938 482406 151174
rect 482170 150618 482406 150854
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 477050 111218 477286 111454
rect 477050 110898 477286 111134
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 471930 57818 472166 58054
rect 471930 57498 472166 57734
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 466810 18098 467046 18334
rect 466810 17778 467046 18014
rect 461690 14378 461926 14614
rect 461690 14058 461926 14294
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 507770 291218 508006 291454
rect 507770 290898 508006 291134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 502650 237818 502886 238054
rect 502650 237498 502886 237734
rect 497530 234098 497766 234334
rect 497530 233778 497766 234014
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 492410 194378 492646 194614
rect 492410 194058 492646 194294
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 487290 154658 487526 154894
rect 487290 154338 487526 154574
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 482170 114938 482406 115174
rect 482170 114618 482406 114854
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 477050 75218 477286 75454
rect 477050 74898 477286 75134
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 471930 21818 472166 22054
rect 471930 21498 472166 21734
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 507770 255218 508006 255454
rect 507770 254898 508006 255134
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 502650 201818 502886 202054
rect 502650 201498 502886 201734
rect 497530 198098 497766 198334
rect 497530 197778 497766 198014
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 492410 158378 492646 158614
rect 492410 158058 492646 158294
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 487290 118658 487526 118894
rect 487290 118338 487526 118574
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 482170 78938 482406 79174
rect 482170 78618 482406 78854
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 477050 39218 477286 39454
rect 477050 38898 477286 39134
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 507770 219218 508006 219454
rect 507770 218898 508006 219134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 502650 165818 502886 166054
rect 502650 165498 502886 165734
rect 497530 162098 497766 162334
rect 497530 161778 497766 162014
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 492410 122378 492646 122614
rect 492410 122058 492646 122294
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 487290 82658 487526 82894
rect 487290 82338 487526 82574
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 482170 42938 482406 43174
rect 482170 42618 482406 42854
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 507770 183218 508006 183454
rect 507770 182898 508006 183134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 502650 129818 502886 130054
rect 502650 129498 502886 129734
rect 497530 126098 497766 126334
rect 497530 125778 497766 126014
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 492410 86378 492646 86614
rect 492410 86058 492646 86294
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 487290 46658 487526 46894
rect 487290 46338 487526 46574
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 482170 6938 482406 7174
rect 482170 6618 482406 6854
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 507770 147218 508006 147454
rect 507770 146898 508006 147134
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 502650 93818 502886 94054
rect 502650 93498 502886 93734
rect 497530 90098 497766 90334
rect 497530 89778 497766 90014
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 492410 50378 492646 50614
rect 492410 50058 492646 50294
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 487290 10658 487526 10894
rect 487290 10338 487526 10574
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 507770 111218 508006 111454
rect 507770 110898 508006 111134
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 502650 57818 502886 58054
rect 502650 57498 502886 57734
rect 497530 54098 497766 54334
rect 497530 53778 497766 54014
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 492410 14378 492646 14614
rect 492410 14058 492646 14294
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 507770 75218 508006 75454
rect 507770 74898 508006 75134
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 502650 21818 502886 22054
rect 502650 21498 502886 21734
rect 497530 18098 497766 18334
rect 497530 17778 497766 18014
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 507770 39218 508006 39454
rect 507770 38898 508006 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 41850 598054
rect 42086 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 72570 598054
rect 72806 597818 103290 598054
rect 103526 597818 134010 598054
rect 134246 597818 164730 598054
rect 164966 597818 195450 598054
rect 195686 597818 226170 598054
rect 226406 597818 256890 598054
rect 257126 597818 287610 598054
rect 287846 597818 318330 598054
rect 318566 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 349050 598054
rect 349286 597818 379770 598054
rect 380006 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 410490 598054
rect 410726 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 441210 598054
rect 441446 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 471930 598054
rect 472166 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 502650 598054
rect 502886 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 41850 597734
rect 42086 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 72570 597734
rect 72806 597498 103290 597734
rect 103526 597498 134010 597734
rect 134246 597498 164730 597734
rect 164966 597498 195450 597734
rect 195686 597498 226170 597734
rect 226406 597498 256890 597734
rect 257126 597498 287610 597734
rect 287846 597498 318330 597734
rect 318566 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 349050 597734
rect 349286 597498 379770 597734
rect 380006 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 410490 597734
rect 410726 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 441210 597734
rect 441446 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 471930 597734
rect 472166 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 502650 597734
rect 502886 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 36730 594334
rect 36966 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 67450 594334
rect 67686 594098 88706 594334
rect 88942 594098 89026 594334
rect 89262 594098 98170 594334
rect 98406 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 128890 594334
rect 129126 594098 159610 594334
rect 159846 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 190330 594334
rect 190566 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 221050 594334
rect 221286 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 251770 594334
rect 252006 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 282490 594334
rect 282726 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 313210 594334
rect 313446 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 343930 594334
rect 344166 594098 374650 594334
rect 374886 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 405370 594334
rect 405606 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 436090 594334
rect 436326 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 466810 594334
rect 467046 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 497530 594334
rect 497766 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 36730 594014
rect 36966 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 67450 594014
rect 67686 593778 88706 594014
rect 88942 593778 89026 594014
rect 89262 593778 98170 594014
rect 98406 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 128890 594014
rect 129126 593778 159610 594014
rect 159846 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 190330 594014
rect 190566 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 221050 594014
rect 221286 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 251770 594014
rect 252006 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 282490 594014
rect 282726 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 313210 594014
rect 313446 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 343930 594014
rect 344166 593778 374650 594014
rect 374886 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 405370 594014
rect 405606 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 436090 594014
rect 436326 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 466810 594014
rect 467046 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 497530 594014
rect 497766 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 31610 590614
rect 31846 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 62330 590614
rect 62566 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 93050 590614
rect 93286 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 123770 590614
rect 124006 590378 154490 590614
rect 154726 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 185210 590614
rect 185446 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 215930 590614
rect 216166 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 246650 590614
rect 246886 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 277370 590614
rect 277606 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 308090 590614
rect 308326 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 338810 590614
rect 339046 590378 369530 590614
rect 369766 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 400250 590614
rect 400486 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 430970 590614
rect 431206 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 461690 590614
rect 461926 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 492410 590614
rect 492646 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 31610 590294
rect 31846 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 62330 590294
rect 62566 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 93050 590294
rect 93286 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 123770 590294
rect 124006 590058 154490 590294
rect 154726 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 185210 590294
rect 185446 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 215930 590294
rect 216166 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 246650 590294
rect 246886 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 277370 590294
rect 277606 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 308090 590294
rect 308326 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 338810 590294
rect 339046 590058 369530 590294
rect 369766 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 400250 590294
rect 400486 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 430970 590294
rect 431206 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 461690 590294
rect 461926 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 492410 590294
rect 492646 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 26490 586894
rect 26726 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 57210 586894
rect 57446 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 87930 586894
rect 88166 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 118650 586894
rect 118886 586658 149370 586894
rect 149606 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 180090 586894
rect 180326 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 210810 586894
rect 211046 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 241530 586894
rect 241766 586658 272250 586894
rect 272486 586658 302970 586894
rect 303206 586658 333690 586894
rect 333926 586658 364410 586894
rect 364646 586658 395130 586894
rect 395366 586658 425850 586894
rect 426086 586658 456570 586894
rect 456806 586658 487290 586894
rect 487526 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 26490 586574
rect 26726 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 57210 586574
rect 57446 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 87930 586574
rect 88166 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 118650 586574
rect 118886 586338 149370 586574
rect 149606 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 180090 586574
rect 180326 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 210810 586574
rect 211046 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 241530 586574
rect 241766 586338 272250 586574
rect 272486 586338 302970 586574
rect 303206 586338 333690 586574
rect 333926 586338 364410 586574
rect 364646 586338 395130 586574
rect 395366 586338 425850 586574
rect 426086 586338 456570 586574
rect 456806 586338 487290 586574
rect 487526 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 21370 583174
rect 21606 582938 52090 583174
rect 52326 582938 82810 583174
rect 83046 582938 113530 583174
rect 113766 582938 144250 583174
rect 144486 582938 174970 583174
rect 175206 582938 205690 583174
rect 205926 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 236410 583174
rect 236646 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 267130 583174
rect 267366 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 297850 583174
rect 298086 582938 328570 583174
rect 328806 582938 359290 583174
rect 359526 582938 390010 583174
rect 390246 582938 420730 583174
rect 420966 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 451450 583174
rect 451686 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 482170 583174
rect 482406 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 21370 582854
rect 21606 582618 52090 582854
rect 52326 582618 82810 582854
rect 83046 582618 113530 582854
rect 113766 582618 144250 582854
rect 144486 582618 174970 582854
rect 175206 582618 205690 582854
rect 205926 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 236410 582854
rect 236646 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 267130 582854
rect 267366 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 297850 582854
rect 298086 582618 328570 582854
rect 328806 582618 359290 582854
rect 359526 582618 390010 582854
rect 390246 582618 420730 582854
rect 420966 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 451450 582854
rect 451686 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 482170 582854
rect 482406 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 16250 579454
rect 16486 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 46970 579454
rect 47206 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 77690 579454
rect 77926 579218 108410 579454
rect 108646 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 139130 579454
rect 139366 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 169850 579454
rect 170086 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 200570 579454
rect 200806 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 231290 579454
rect 231526 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 262010 579454
rect 262246 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 292730 579454
rect 292966 579218 323450 579454
rect 323686 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 354170 579454
rect 354406 579218 384890 579454
rect 385126 579218 415610 579454
rect 415846 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 446330 579454
rect 446566 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 477050 579454
rect 477286 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 507770 579454
rect 508006 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 16250 579134
rect 16486 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 46970 579134
rect 47206 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 77690 579134
rect 77926 578898 108410 579134
rect 108646 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 139130 579134
rect 139366 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 169850 579134
rect 170086 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 200570 579134
rect 200806 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 231290 579134
rect 231526 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 262010 579134
rect 262246 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 292730 579134
rect 292966 578898 323450 579134
rect 323686 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 354170 579134
rect 354406 578898 384890 579134
rect 385126 578898 415610 579134
rect 415846 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 446330 579134
rect 446566 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 477050 579134
rect 477286 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 507770 579134
rect 508006 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 41850 562054
rect 42086 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 72570 562054
rect 72806 561818 103290 562054
rect 103526 561818 134010 562054
rect 134246 561818 164730 562054
rect 164966 561818 195450 562054
rect 195686 561818 226170 562054
rect 226406 561818 256890 562054
rect 257126 561818 287610 562054
rect 287846 561818 318330 562054
rect 318566 561818 349050 562054
rect 349286 561818 379770 562054
rect 380006 561818 410490 562054
rect 410726 561818 441210 562054
rect 441446 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 471930 562054
rect 472166 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 502650 562054
rect 502886 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 41850 561734
rect 42086 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 72570 561734
rect 72806 561498 103290 561734
rect 103526 561498 134010 561734
rect 134246 561498 164730 561734
rect 164966 561498 195450 561734
rect 195686 561498 226170 561734
rect 226406 561498 256890 561734
rect 257126 561498 287610 561734
rect 287846 561498 318330 561734
rect 318566 561498 349050 561734
rect 349286 561498 379770 561734
rect 380006 561498 410490 561734
rect 410726 561498 441210 561734
rect 441446 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 471930 561734
rect 472166 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 502650 561734
rect 502886 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 36730 558334
rect 36966 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 67450 558334
rect 67686 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 98170 558334
rect 98406 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 128890 558334
rect 129126 558098 159610 558334
rect 159846 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 190330 558334
rect 190566 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 221050 558334
rect 221286 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 251770 558334
rect 252006 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 282490 558334
rect 282726 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 313210 558334
rect 313446 558098 343930 558334
rect 344166 558098 374650 558334
rect 374886 558098 405370 558334
rect 405606 558098 436090 558334
rect 436326 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 466810 558334
rect 467046 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 497530 558334
rect 497766 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 36730 558014
rect 36966 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 67450 558014
rect 67686 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 98170 558014
rect 98406 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 128890 558014
rect 129126 557778 159610 558014
rect 159846 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 190330 558014
rect 190566 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 221050 558014
rect 221286 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 251770 558014
rect 252006 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 282490 558014
rect 282726 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 313210 558014
rect 313446 557778 343930 558014
rect 344166 557778 374650 558014
rect 374886 557778 405370 558014
rect 405606 557778 436090 558014
rect 436326 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 466810 558014
rect 467046 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 497530 558014
rect 497766 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 31610 554614
rect 31846 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 62330 554614
rect 62566 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 93050 554614
rect 93286 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 123770 554614
rect 124006 554378 154490 554614
rect 154726 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 185210 554614
rect 185446 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 215930 554614
rect 216166 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 246650 554614
rect 246886 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 277370 554614
rect 277606 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 308090 554614
rect 308326 554378 338810 554614
rect 339046 554378 369530 554614
rect 369766 554378 400250 554614
rect 400486 554378 430970 554614
rect 431206 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 461690 554614
rect 461926 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 492410 554614
rect 492646 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 31610 554294
rect 31846 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 62330 554294
rect 62566 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 93050 554294
rect 93286 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 123770 554294
rect 124006 554058 154490 554294
rect 154726 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 185210 554294
rect 185446 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 215930 554294
rect 216166 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 246650 554294
rect 246886 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 277370 554294
rect 277606 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 308090 554294
rect 308326 554058 338810 554294
rect 339046 554058 369530 554294
rect 369766 554058 400250 554294
rect 400486 554058 430970 554294
rect 431206 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 461690 554294
rect 461926 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 492410 554294
rect 492646 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 26490 550894
rect 26726 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 57210 550894
rect 57446 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 87930 550894
rect 88166 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 118650 550894
rect 118886 550658 149370 550894
rect 149606 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 180090 550894
rect 180326 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 210810 550894
rect 211046 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 241530 550894
rect 241766 550658 272250 550894
rect 272486 550658 302970 550894
rect 303206 550658 333690 550894
rect 333926 550658 364410 550894
rect 364646 550658 395130 550894
rect 395366 550658 425850 550894
rect 426086 550658 456570 550894
rect 456806 550658 487290 550894
rect 487526 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 26490 550574
rect 26726 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 57210 550574
rect 57446 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 87930 550574
rect 88166 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 118650 550574
rect 118886 550338 149370 550574
rect 149606 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 180090 550574
rect 180326 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 210810 550574
rect 211046 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 241530 550574
rect 241766 550338 272250 550574
rect 272486 550338 302970 550574
rect 303206 550338 333690 550574
rect 333926 550338 364410 550574
rect 364646 550338 395130 550574
rect 395366 550338 425850 550574
rect 426086 550338 456570 550574
rect 456806 550338 487290 550574
rect 487526 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 21370 547174
rect 21606 546938 52090 547174
rect 52326 546938 82810 547174
rect 83046 546938 113530 547174
rect 113766 546938 144250 547174
rect 144486 546938 174970 547174
rect 175206 546938 205690 547174
rect 205926 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 236410 547174
rect 236646 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 267130 547174
rect 267366 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 297850 547174
rect 298086 546938 328570 547174
rect 328806 546938 359290 547174
rect 359526 546938 390010 547174
rect 390246 546938 420730 547174
rect 420966 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 451450 547174
rect 451686 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 482170 547174
rect 482406 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 21370 546854
rect 21606 546618 52090 546854
rect 52326 546618 82810 546854
rect 83046 546618 113530 546854
rect 113766 546618 144250 546854
rect 144486 546618 174970 546854
rect 175206 546618 205690 546854
rect 205926 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 236410 546854
rect 236646 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 267130 546854
rect 267366 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 297850 546854
rect 298086 546618 328570 546854
rect 328806 546618 359290 546854
rect 359526 546618 390010 546854
rect 390246 546618 420730 546854
rect 420966 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 451450 546854
rect 451686 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 482170 546854
rect 482406 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 16250 543454
rect 16486 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 46970 543454
rect 47206 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 77690 543454
rect 77926 543218 108410 543454
rect 108646 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 139130 543454
rect 139366 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 169850 543454
rect 170086 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 200570 543454
rect 200806 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 231290 543454
rect 231526 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 262010 543454
rect 262246 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 292730 543454
rect 292966 543218 323450 543454
rect 323686 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 354170 543454
rect 354406 543218 384890 543454
rect 385126 543218 415610 543454
rect 415846 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 446330 543454
rect 446566 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 477050 543454
rect 477286 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 507770 543454
rect 508006 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 16250 543134
rect 16486 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 46970 543134
rect 47206 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 77690 543134
rect 77926 542898 108410 543134
rect 108646 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 139130 543134
rect 139366 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 169850 543134
rect 170086 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 200570 543134
rect 200806 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 231290 543134
rect 231526 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 262010 543134
rect 262246 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 292730 543134
rect 292966 542898 323450 543134
rect 323686 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 354170 543134
rect 354406 542898 384890 543134
rect 385126 542898 415610 543134
rect 415846 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 446330 543134
rect 446566 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 477050 543134
rect 477286 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 507770 543134
rect 508006 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 41850 526054
rect 42086 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 72570 526054
rect 72806 525818 103290 526054
rect 103526 525818 134010 526054
rect 134246 525818 164730 526054
rect 164966 525818 195450 526054
rect 195686 525818 226170 526054
rect 226406 525818 256890 526054
rect 257126 525818 287610 526054
rect 287846 525818 318330 526054
rect 318566 525818 349050 526054
rect 349286 525818 379770 526054
rect 380006 525818 410490 526054
rect 410726 525818 441210 526054
rect 441446 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 471930 526054
rect 472166 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 502650 526054
rect 502886 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 41850 525734
rect 42086 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 72570 525734
rect 72806 525498 103290 525734
rect 103526 525498 134010 525734
rect 134246 525498 164730 525734
rect 164966 525498 195450 525734
rect 195686 525498 226170 525734
rect 226406 525498 256890 525734
rect 257126 525498 287610 525734
rect 287846 525498 318330 525734
rect 318566 525498 349050 525734
rect 349286 525498 379770 525734
rect 380006 525498 410490 525734
rect 410726 525498 441210 525734
rect 441446 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 471930 525734
rect 472166 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 502650 525734
rect 502886 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 36730 522334
rect 36966 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 67450 522334
rect 67686 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 98170 522334
rect 98406 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 128890 522334
rect 129126 522098 159610 522334
rect 159846 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 190330 522334
rect 190566 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 221050 522334
rect 221286 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 251770 522334
rect 252006 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 282490 522334
rect 282726 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 313210 522334
rect 313446 522098 343930 522334
rect 344166 522098 374650 522334
rect 374886 522098 405370 522334
rect 405606 522098 436090 522334
rect 436326 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 466810 522334
rect 467046 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 497530 522334
rect 497766 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 36730 522014
rect 36966 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 67450 522014
rect 67686 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 98170 522014
rect 98406 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 128890 522014
rect 129126 521778 159610 522014
rect 159846 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 190330 522014
rect 190566 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 221050 522014
rect 221286 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 251770 522014
rect 252006 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 282490 522014
rect 282726 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 313210 522014
rect 313446 521778 343930 522014
rect 344166 521778 374650 522014
rect 374886 521778 405370 522014
rect 405606 521778 436090 522014
rect 436326 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 466810 522014
rect 467046 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 497530 522014
rect 497766 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 31610 518614
rect 31846 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 62330 518614
rect 62566 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 93050 518614
rect 93286 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 123770 518614
rect 124006 518378 154490 518614
rect 154726 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 185210 518614
rect 185446 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 215930 518614
rect 216166 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 246650 518614
rect 246886 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 277370 518614
rect 277606 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 308090 518614
rect 308326 518378 338810 518614
rect 339046 518378 369530 518614
rect 369766 518378 400250 518614
rect 400486 518378 430970 518614
rect 431206 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 461690 518614
rect 461926 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 492410 518614
rect 492646 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 31610 518294
rect 31846 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 62330 518294
rect 62566 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 93050 518294
rect 93286 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 123770 518294
rect 124006 518058 154490 518294
rect 154726 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 185210 518294
rect 185446 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 215930 518294
rect 216166 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 246650 518294
rect 246886 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 277370 518294
rect 277606 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 308090 518294
rect 308326 518058 338810 518294
rect 339046 518058 369530 518294
rect 369766 518058 400250 518294
rect 400486 518058 430970 518294
rect 431206 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 461690 518294
rect 461926 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 492410 518294
rect 492646 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 26490 514894
rect 26726 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 57210 514894
rect 57446 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 87930 514894
rect 88166 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 118650 514894
rect 118886 514658 149370 514894
rect 149606 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 180090 514894
rect 180326 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 210810 514894
rect 211046 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 241530 514894
rect 241766 514658 272250 514894
rect 272486 514658 302970 514894
rect 303206 514658 333690 514894
rect 333926 514658 364410 514894
rect 364646 514658 395130 514894
rect 395366 514658 425850 514894
rect 426086 514658 456570 514894
rect 456806 514658 487290 514894
rect 487526 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 26490 514574
rect 26726 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 57210 514574
rect 57446 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 87930 514574
rect 88166 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 118650 514574
rect 118886 514338 149370 514574
rect 149606 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 180090 514574
rect 180326 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 210810 514574
rect 211046 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 241530 514574
rect 241766 514338 272250 514574
rect 272486 514338 302970 514574
rect 303206 514338 333690 514574
rect 333926 514338 364410 514574
rect 364646 514338 395130 514574
rect 395366 514338 425850 514574
rect 426086 514338 456570 514574
rect 456806 514338 487290 514574
rect 487526 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 21370 511174
rect 21606 510938 52090 511174
rect 52326 510938 82810 511174
rect 83046 510938 113530 511174
rect 113766 510938 144250 511174
rect 144486 510938 174970 511174
rect 175206 510938 205690 511174
rect 205926 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 236410 511174
rect 236646 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 267130 511174
rect 267366 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 297850 511174
rect 298086 510938 328570 511174
rect 328806 510938 359290 511174
rect 359526 510938 390010 511174
rect 390246 510938 420730 511174
rect 420966 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 451450 511174
rect 451686 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 482170 511174
rect 482406 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 21370 510854
rect 21606 510618 52090 510854
rect 52326 510618 82810 510854
rect 83046 510618 113530 510854
rect 113766 510618 144250 510854
rect 144486 510618 174970 510854
rect 175206 510618 205690 510854
rect 205926 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 236410 510854
rect 236646 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 267130 510854
rect 267366 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 297850 510854
rect 298086 510618 328570 510854
rect 328806 510618 359290 510854
rect 359526 510618 390010 510854
rect 390246 510618 420730 510854
rect 420966 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 451450 510854
rect 451686 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 482170 510854
rect 482406 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 16250 507454
rect 16486 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 46970 507454
rect 47206 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 77690 507454
rect 77926 507218 108410 507454
rect 108646 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 139130 507454
rect 139366 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 169850 507454
rect 170086 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 200570 507454
rect 200806 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 231290 507454
rect 231526 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 262010 507454
rect 262246 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 292730 507454
rect 292966 507218 323450 507454
rect 323686 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 354170 507454
rect 354406 507218 384890 507454
rect 385126 507218 415610 507454
rect 415846 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 446330 507454
rect 446566 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 477050 507454
rect 477286 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 507770 507454
rect 508006 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 16250 507134
rect 16486 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 46970 507134
rect 47206 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 77690 507134
rect 77926 506898 108410 507134
rect 108646 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 139130 507134
rect 139366 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 169850 507134
rect 170086 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 200570 507134
rect 200806 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 231290 507134
rect 231526 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 262010 507134
rect 262246 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 292730 507134
rect 292966 506898 323450 507134
rect 323686 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 354170 507134
rect 354406 506898 384890 507134
rect 385126 506898 415610 507134
rect 415846 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 446330 507134
rect 446566 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 477050 507134
rect 477286 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 507770 507134
rect 508006 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 41850 490054
rect 42086 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 72570 490054
rect 72806 489818 103290 490054
rect 103526 489818 134010 490054
rect 134246 489818 164730 490054
rect 164966 489818 195450 490054
rect 195686 489818 226170 490054
rect 226406 489818 256890 490054
rect 257126 489818 287610 490054
rect 287846 489818 318330 490054
rect 318566 489818 349050 490054
rect 349286 489818 379770 490054
rect 380006 489818 410490 490054
rect 410726 489818 441210 490054
rect 441446 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 471930 490054
rect 472166 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 502650 490054
rect 502886 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 41850 489734
rect 42086 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 72570 489734
rect 72806 489498 103290 489734
rect 103526 489498 134010 489734
rect 134246 489498 164730 489734
rect 164966 489498 195450 489734
rect 195686 489498 226170 489734
rect 226406 489498 256890 489734
rect 257126 489498 287610 489734
rect 287846 489498 318330 489734
rect 318566 489498 349050 489734
rect 349286 489498 379770 489734
rect 380006 489498 410490 489734
rect 410726 489498 441210 489734
rect 441446 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 471930 489734
rect 472166 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 502650 489734
rect 502886 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 36730 486334
rect 36966 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 67450 486334
rect 67686 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 98170 486334
rect 98406 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 128890 486334
rect 129126 486098 159610 486334
rect 159846 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 190330 486334
rect 190566 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 221050 486334
rect 221286 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 251770 486334
rect 252006 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 282490 486334
rect 282726 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 313210 486334
rect 313446 486098 343930 486334
rect 344166 486098 374650 486334
rect 374886 486098 405370 486334
rect 405606 486098 436090 486334
rect 436326 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 466810 486334
rect 467046 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 497530 486334
rect 497766 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 36730 486014
rect 36966 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 67450 486014
rect 67686 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 98170 486014
rect 98406 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 128890 486014
rect 129126 485778 159610 486014
rect 159846 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 190330 486014
rect 190566 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 221050 486014
rect 221286 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 251770 486014
rect 252006 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 282490 486014
rect 282726 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 313210 486014
rect 313446 485778 343930 486014
rect 344166 485778 374650 486014
rect 374886 485778 405370 486014
rect 405606 485778 436090 486014
rect 436326 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 466810 486014
rect 467046 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 497530 486014
rect 497766 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 31610 482614
rect 31846 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 62330 482614
rect 62566 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 93050 482614
rect 93286 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 123770 482614
rect 124006 482378 154490 482614
rect 154726 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 185210 482614
rect 185446 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 215930 482614
rect 216166 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 246650 482614
rect 246886 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 277370 482614
rect 277606 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 308090 482614
rect 308326 482378 338810 482614
rect 339046 482378 369530 482614
rect 369766 482378 400250 482614
rect 400486 482378 430970 482614
rect 431206 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 461690 482614
rect 461926 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 492410 482614
rect 492646 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 31610 482294
rect 31846 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 62330 482294
rect 62566 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 93050 482294
rect 93286 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 123770 482294
rect 124006 482058 154490 482294
rect 154726 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 185210 482294
rect 185446 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 215930 482294
rect 216166 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 246650 482294
rect 246886 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 277370 482294
rect 277606 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 308090 482294
rect 308326 482058 338810 482294
rect 339046 482058 369530 482294
rect 369766 482058 400250 482294
rect 400486 482058 430970 482294
rect 431206 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 461690 482294
rect 461926 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 492410 482294
rect 492646 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 26490 478894
rect 26726 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 57210 478894
rect 57446 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 87930 478894
rect 88166 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 118650 478894
rect 118886 478658 149370 478894
rect 149606 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 180090 478894
rect 180326 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 210810 478894
rect 211046 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 241530 478894
rect 241766 478658 272250 478894
rect 272486 478658 302970 478894
rect 303206 478658 333690 478894
rect 333926 478658 364410 478894
rect 364646 478658 395130 478894
rect 395366 478658 425850 478894
rect 426086 478658 456570 478894
rect 456806 478658 487290 478894
rect 487526 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 26490 478574
rect 26726 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 57210 478574
rect 57446 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 87930 478574
rect 88166 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 118650 478574
rect 118886 478338 149370 478574
rect 149606 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 180090 478574
rect 180326 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 210810 478574
rect 211046 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 241530 478574
rect 241766 478338 272250 478574
rect 272486 478338 302970 478574
rect 303206 478338 333690 478574
rect 333926 478338 364410 478574
rect 364646 478338 395130 478574
rect 395366 478338 425850 478574
rect 426086 478338 456570 478574
rect 456806 478338 487290 478574
rect 487526 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 21370 475174
rect 21606 474938 52090 475174
rect 52326 474938 82810 475174
rect 83046 474938 113530 475174
rect 113766 474938 144250 475174
rect 144486 474938 174970 475174
rect 175206 474938 205690 475174
rect 205926 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 236410 475174
rect 236646 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 267130 475174
rect 267366 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 297850 475174
rect 298086 474938 328570 475174
rect 328806 474938 359290 475174
rect 359526 474938 390010 475174
rect 390246 474938 420730 475174
rect 420966 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 451450 475174
rect 451686 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 482170 475174
rect 482406 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 21370 474854
rect 21606 474618 52090 474854
rect 52326 474618 82810 474854
rect 83046 474618 113530 474854
rect 113766 474618 144250 474854
rect 144486 474618 174970 474854
rect 175206 474618 205690 474854
rect 205926 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 236410 474854
rect 236646 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 267130 474854
rect 267366 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 297850 474854
rect 298086 474618 328570 474854
rect 328806 474618 359290 474854
rect 359526 474618 390010 474854
rect 390246 474618 420730 474854
rect 420966 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 451450 474854
rect 451686 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 482170 474854
rect 482406 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 16250 471454
rect 16486 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 46970 471454
rect 47206 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 77690 471454
rect 77926 471218 108410 471454
rect 108646 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 139130 471454
rect 139366 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 169850 471454
rect 170086 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 200570 471454
rect 200806 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 231290 471454
rect 231526 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 262010 471454
rect 262246 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 292730 471454
rect 292966 471218 323450 471454
rect 323686 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 354170 471454
rect 354406 471218 384890 471454
rect 385126 471218 415610 471454
rect 415846 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 446330 471454
rect 446566 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 477050 471454
rect 477286 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 507770 471454
rect 508006 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 16250 471134
rect 16486 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 46970 471134
rect 47206 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 77690 471134
rect 77926 470898 108410 471134
rect 108646 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 139130 471134
rect 139366 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 169850 471134
rect 170086 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 200570 471134
rect 200806 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 231290 471134
rect 231526 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 262010 471134
rect 262246 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 292730 471134
rect 292966 470898 323450 471134
rect 323686 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 354170 471134
rect 354406 470898 384890 471134
rect 385126 470898 415610 471134
rect 415846 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 446330 471134
rect 446566 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 477050 471134
rect 477286 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 507770 471134
rect 508006 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 41850 454054
rect 42086 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 72570 454054
rect 72806 453818 103290 454054
rect 103526 453818 134010 454054
rect 134246 453818 164730 454054
rect 164966 453818 195450 454054
rect 195686 453818 226170 454054
rect 226406 453818 256890 454054
rect 257126 453818 287610 454054
rect 287846 453818 318330 454054
rect 318566 453818 349050 454054
rect 349286 453818 379770 454054
rect 380006 453818 410490 454054
rect 410726 453818 441210 454054
rect 441446 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 471930 454054
rect 472166 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 502650 454054
rect 502886 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 41850 453734
rect 42086 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 72570 453734
rect 72806 453498 103290 453734
rect 103526 453498 134010 453734
rect 134246 453498 164730 453734
rect 164966 453498 195450 453734
rect 195686 453498 226170 453734
rect 226406 453498 256890 453734
rect 257126 453498 287610 453734
rect 287846 453498 318330 453734
rect 318566 453498 349050 453734
rect 349286 453498 379770 453734
rect 380006 453498 410490 453734
rect 410726 453498 441210 453734
rect 441446 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 471930 453734
rect 472166 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 502650 453734
rect 502886 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 36730 450334
rect 36966 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 67450 450334
rect 67686 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 98170 450334
rect 98406 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 128890 450334
rect 129126 450098 159610 450334
rect 159846 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 190330 450334
rect 190566 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 221050 450334
rect 221286 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 251770 450334
rect 252006 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 282490 450334
rect 282726 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 313210 450334
rect 313446 450098 343930 450334
rect 344166 450098 374650 450334
rect 374886 450098 405370 450334
rect 405606 450098 436090 450334
rect 436326 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 466810 450334
rect 467046 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 497530 450334
rect 497766 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 36730 450014
rect 36966 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 67450 450014
rect 67686 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 98170 450014
rect 98406 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 128890 450014
rect 129126 449778 159610 450014
rect 159846 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 190330 450014
rect 190566 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 221050 450014
rect 221286 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 251770 450014
rect 252006 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 282490 450014
rect 282726 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 313210 450014
rect 313446 449778 343930 450014
rect 344166 449778 374650 450014
rect 374886 449778 405370 450014
rect 405606 449778 436090 450014
rect 436326 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 466810 450014
rect 467046 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 497530 450014
rect 497766 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 31610 446614
rect 31846 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 62330 446614
rect 62566 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 93050 446614
rect 93286 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 123770 446614
rect 124006 446378 154490 446614
rect 154726 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 185210 446614
rect 185446 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 215930 446614
rect 216166 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 246650 446614
rect 246886 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 277370 446614
rect 277606 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 308090 446614
rect 308326 446378 338810 446614
rect 339046 446378 369530 446614
rect 369766 446378 400250 446614
rect 400486 446378 430970 446614
rect 431206 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 461690 446614
rect 461926 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 492410 446614
rect 492646 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 31610 446294
rect 31846 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 62330 446294
rect 62566 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 93050 446294
rect 93286 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 123770 446294
rect 124006 446058 154490 446294
rect 154726 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 185210 446294
rect 185446 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 215930 446294
rect 216166 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 246650 446294
rect 246886 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 277370 446294
rect 277606 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 308090 446294
rect 308326 446058 338810 446294
rect 339046 446058 369530 446294
rect 369766 446058 400250 446294
rect 400486 446058 430970 446294
rect 431206 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 461690 446294
rect 461926 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 492410 446294
rect 492646 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 26490 442894
rect 26726 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 57210 442894
rect 57446 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 87930 442894
rect 88166 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 118650 442894
rect 118886 442658 149370 442894
rect 149606 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 180090 442894
rect 180326 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 210810 442894
rect 211046 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 241530 442894
rect 241766 442658 272250 442894
rect 272486 442658 302970 442894
rect 303206 442658 333690 442894
rect 333926 442658 364410 442894
rect 364646 442658 395130 442894
rect 395366 442658 425850 442894
rect 426086 442658 456570 442894
rect 456806 442658 487290 442894
rect 487526 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 26490 442574
rect 26726 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 57210 442574
rect 57446 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 87930 442574
rect 88166 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 118650 442574
rect 118886 442338 149370 442574
rect 149606 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 180090 442574
rect 180326 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 210810 442574
rect 211046 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 241530 442574
rect 241766 442338 272250 442574
rect 272486 442338 302970 442574
rect 303206 442338 333690 442574
rect 333926 442338 364410 442574
rect 364646 442338 395130 442574
rect 395366 442338 425850 442574
rect 426086 442338 456570 442574
rect 456806 442338 487290 442574
rect 487526 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 21370 439174
rect 21606 438938 52090 439174
rect 52326 438938 82810 439174
rect 83046 438938 113530 439174
rect 113766 438938 144250 439174
rect 144486 438938 174970 439174
rect 175206 438938 205690 439174
rect 205926 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 236410 439174
rect 236646 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 267130 439174
rect 267366 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 297850 439174
rect 298086 438938 328570 439174
rect 328806 438938 359290 439174
rect 359526 438938 390010 439174
rect 390246 438938 420730 439174
rect 420966 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 451450 439174
rect 451686 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 482170 439174
rect 482406 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 21370 438854
rect 21606 438618 52090 438854
rect 52326 438618 82810 438854
rect 83046 438618 113530 438854
rect 113766 438618 144250 438854
rect 144486 438618 174970 438854
rect 175206 438618 205690 438854
rect 205926 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 236410 438854
rect 236646 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 267130 438854
rect 267366 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 297850 438854
rect 298086 438618 328570 438854
rect 328806 438618 359290 438854
rect 359526 438618 390010 438854
rect 390246 438618 420730 438854
rect 420966 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 451450 438854
rect 451686 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 482170 438854
rect 482406 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 16250 435454
rect 16486 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 46970 435454
rect 47206 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 77690 435454
rect 77926 435218 108410 435454
rect 108646 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 139130 435454
rect 139366 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 169850 435454
rect 170086 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 200570 435454
rect 200806 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 231290 435454
rect 231526 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 262010 435454
rect 262246 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 292730 435454
rect 292966 435218 323450 435454
rect 323686 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 354170 435454
rect 354406 435218 384890 435454
rect 385126 435218 415610 435454
rect 415846 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 446330 435454
rect 446566 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 477050 435454
rect 477286 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 507770 435454
rect 508006 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 16250 435134
rect 16486 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 46970 435134
rect 47206 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 77690 435134
rect 77926 434898 108410 435134
rect 108646 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 139130 435134
rect 139366 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 169850 435134
rect 170086 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 200570 435134
rect 200806 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 231290 435134
rect 231526 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 262010 435134
rect 262246 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 292730 435134
rect 292966 434898 323450 435134
rect 323686 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 354170 435134
rect 354406 434898 384890 435134
rect 385126 434898 415610 435134
rect 415846 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 446330 435134
rect 446566 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 477050 435134
rect 477286 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 507770 435134
rect 508006 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 41850 418054
rect 42086 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 72570 418054
rect 72806 417818 103290 418054
rect 103526 417818 134010 418054
rect 134246 417818 164730 418054
rect 164966 417818 195450 418054
rect 195686 417818 226170 418054
rect 226406 417818 256890 418054
rect 257126 417818 287610 418054
rect 287846 417818 318330 418054
rect 318566 417818 349050 418054
rect 349286 417818 379770 418054
rect 380006 417818 410490 418054
rect 410726 417818 441210 418054
rect 441446 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 471930 418054
rect 472166 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 502650 418054
rect 502886 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 41850 417734
rect 42086 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 72570 417734
rect 72806 417498 103290 417734
rect 103526 417498 134010 417734
rect 134246 417498 164730 417734
rect 164966 417498 195450 417734
rect 195686 417498 226170 417734
rect 226406 417498 256890 417734
rect 257126 417498 287610 417734
rect 287846 417498 318330 417734
rect 318566 417498 349050 417734
rect 349286 417498 379770 417734
rect 380006 417498 410490 417734
rect 410726 417498 441210 417734
rect 441446 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 471930 417734
rect 472166 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 502650 417734
rect 502886 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 36730 414334
rect 36966 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 67450 414334
rect 67686 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 98170 414334
rect 98406 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 128890 414334
rect 129126 414098 159610 414334
rect 159846 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 190330 414334
rect 190566 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 221050 414334
rect 221286 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 251770 414334
rect 252006 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 282490 414334
rect 282726 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 313210 414334
rect 313446 414098 343930 414334
rect 344166 414098 374650 414334
rect 374886 414098 405370 414334
rect 405606 414098 436090 414334
rect 436326 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 466810 414334
rect 467046 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 497530 414334
rect 497766 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 36730 414014
rect 36966 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 67450 414014
rect 67686 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 98170 414014
rect 98406 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 128890 414014
rect 129126 413778 159610 414014
rect 159846 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 190330 414014
rect 190566 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 221050 414014
rect 221286 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 251770 414014
rect 252006 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 282490 414014
rect 282726 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 313210 414014
rect 313446 413778 343930 414014
rect 344166 413778 374650 414014
rect 374886 413778 405370 414014
rect 405606 413778 436090 414014
rect 436326 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 466810 414014
rect 467046 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 497530 414014
rect 497766 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 31610 410614
rect 31846 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 62330 410614
rect 62566 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 93050 410614
rect 93286 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 123770 410614
rect 124006 410378 154490 410614
rect 154726 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 185210 410614
rect 185446 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 215930 410614
rect 216166 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 246650 410614
rect 246886 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 277370 410614
rect 277606 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 308090 410614
rect 308326 410378 338810 410614
rect 339046 410378 369530 410614
rect 369766 410378 400250 410614
rect 400486 410378 430970 410614
rect 431206 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 461690 410614
rect 461926 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 492410 410614
rect 492646 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 31610 410294
rect 31846 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 62330 410294
rect 62566 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 93050 410294
rect 93286 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 123770 410294
rect 124006 410058 154490 410294
rect 154726 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 185210 410294
rect 185446 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 215930 410294
rect 216166 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 246650 410294
rect 246886 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 277370 410294
rect 277606 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 308090 410294
rect 308326 410058 338810 410294
rect 339046 410058 369530 410294
rect 369766 410058 400250 410294
rect 400486 410058 430970 410294
rect 431206 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 461690 410294
rect 461926 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 492410 410294
rect 492646 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 26490 406894
rect 26726 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 57210 406894
rect 57446 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 87930 406894
rect 88166 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 118650 406894
rect 118886 406658 149370 406894
rect 149606 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 180090 406894
rect 180326 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 210810 406894
rect 211046 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 241530 406894
rect 241766 406658 272250 406894
rect 272486 406658 302970 406894
rect 303206 406658 333690 406894
rect 333926 406658 364410 406894
rect 364646 406658 395130 406894
rect 395366 406658 425850 406894
rect 426086 406658 456570 406894
rect 456806 406658 487290 406894
rect 487526 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 26490 406574
rect 26726 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 57210 406574
rect 57446 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 87930 406574
rect 88166 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 118650 406574
rect 118886 406338 149370 406574
rect 149606 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 180090 406574
rect 180326 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 210810 406574
rect 211046 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 241530 406574
rect 241766 406338 272250 406574
rect 272486 406338 302970 406574
rect 303206 406338 333690 406574
rect 333926 406338 364410 406574
rect 364646 406338 395130 406574
rect 395366 406338 425850 406574
rect 426086 406338 456570 406574
rect 456806 406338 487290 406574
rect 487526 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 21370 403174
rect 21606 402938 52090 403174
rect 52326 402938 82810 403174
rect 83046 402938 113530 403174
rect 113766 402938 144250 403174
rect 144486 402938 174970 403174
rect 175206 402938 205690 403174
rect 205926 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 236410 403174
rect 236646 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 267130 403174
rect 267366 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 297850 403174
rect 298086 402938 328570 403174
rect 328806 402938 359290 403174
rect 359526 402938 390010 403174
rect 390246 402938 420730 403174
rect 420966 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 451450 403174
rect 451686 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 482170 403174
rect 482406 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 21370 402854
rect 21606 402618 52090 402854
rect 52326 402618 82810 402854
rect 83046 402618 113530 402854
rect 113766 402618 144250 402854
rect 144486 402618 174970 402854
rect 175206 402618 205690 402854
rect 205926 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 236410 402854
rect 236646 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 267130 402854
rect 267366 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 297850 402854
rect 298086 402618 328570 402854
rect 328806 402618 359290 402854
rect 359526 402618 390010 402854
rect 390246 402618 420730 402854
rect 420966 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 451450 402854
rect 451686 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 482170 402854
rect 482406 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 16250 399454
rect 16486 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 46970 399454
rect 47206 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 77690 399454
rect 77926 399218 108410 399454
rect 108646 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 139130 399454
rect 139366 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 169850 399454
rect 170086 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 200570 399454
rect 200806 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 231290 399454
rect 231526 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 262010 399454
rect 262246 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 292730 399454
rect 292966 399218 323450 399454
rect 323686 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 354170 399454
rect 354406 399218 384890 399454
rect 385126 399218 415610 399454
rect 415846 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 446330 399454
rect 446566 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 477050 399454
rect 477286 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 507770 399454
rect 508006 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 16250 399134
rect 16486 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 46970 399134
rect 47206 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 77690 399134
rect 77926 398898 108410 399134
rect 108646 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 139130 399134
rect 139366 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 169850 399134
rect 170086 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 200570 399134
rect 200806 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 231290 399134
rect 231526 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 262010 399134
rect 262246 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 292730 399134
rect 292966 398898 323450 399134
rect 323686 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 354170 399134
rect 354406 398898 384890 399134
rect 385126 398898 415610 399134
rect 415846 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 446330 399134
rect 446566 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 477050 399134
rect 477286 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 507770 399134
rect 508006 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 41850 382054
rect 42086 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 72570 382054
rect 72806 381818 103290 382054
rect 103526 381818 134010 382054
rect 134246 381818 164730 382054
rect 164966 381818 195450 382054
rect 195686 381818 226170 382054
rect 226406 381818 256890 382054
rect 257126 381818 287610 382054
rect 287846 381818 318330 382054
rect 318566 381818 349050 382054
rect 349286 381818 379770 382054
rect 380006 381818 410490 382054
rect 410726 381818 441210 382054
rect 441446 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 471930 382054
rect 472166 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 502650 382054
rect 502886 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 41850 381734
rect 42086 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 72570 381734
rect 72806 381498 103290 381734
rect 103526 381498 134010 381734
rect 134246 381498 164730 381734
rect 164966 381498 195450 381734
rect 195686 381498 226170 381734
rect 226406 381498 256890 381734
rect 257126 381498 287610 381734
rect 287846 381498 318330 381734
rect 318566 381498 349050 381734
rect 349286 381498 379770 381734
rect 380006 381498 410490 381734
rect 410726 381498 441210 381734
rect 441446 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 471930 381734
rect 472166 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 502650 381734
rect 502886 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 36730 378334
rect 36966 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 67450 378334
rect 67686 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 98170 378334
rect 98406 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 128890 378334
rect 129126 378098 159610 378334
rect 159846 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 190330 378334
rect 190566 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 221050 378334
rect 221286 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 251770 378334
rect 252006 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 282490 378334
rect 282726 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 313210 378334
rect 313446 378098 343930 378334
rect 344166 378098 374650 378334
rect 374886 378098 405370 378334
rect 405606 378098 436090 378334
rect 436326 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 466810 378334
rect 467046 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 497530 378334
rect 497766 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 36730 378014
rect 36966 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 67450 378014
rect 67686 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 98170 378014
rect 98406 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 128890 378014
rect 129126 377778 159610 378014
rect 159846 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 190330 378014
rect 190566 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 221050 378014
rect 221286 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 251770 378014
rect 252006 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 282490 378014
rect 282726 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 313210 378014
rect 313446 377778 343930 378014
rect 344166 377778 374650 378014
rect 374886 377778 405370 378014
rect 405606 377778 436090 378014
rect 436326 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 466810 378014
rect 467046 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 497530 378014
rect 497766 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 31610 374614
rect 31846 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 62330 374614
rect 62566 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 93050 374614
rect 93286 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 123770 374614
rect 124006 374378 154490 374614
rect 154726 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 185210 374614
rect 185446 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 215930 374614
rect 216166 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 246650 374614
rect 246886 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 277370 374614
rect 277606 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 308090 374614
rect 308326 374378 338810 374614
rect 339046 374378 369530 374614
rect 369766 374378 400250 374614
rect 400486 374378 430970 374614
rect 431206 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 461690 374614
rect 461926 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 492410 374614
rect 492646 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 31610 374294
rect 31846 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 62330 374294
rect 62566 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 93050 374294
rect 93286 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 123770 374294
rect 124006 374058 154490 374294
rect 154726 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 185210 374294
rect 185446 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 215930 374294
rect 216166 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 246650 374294
rect 246886 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 277370 374294
rect 277606 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 308090 374294
rect 308326 374058 338810 374294
rect 339046 374058 369530 374294
rect 369766 374058 400250 374294
rect 400486 374058 430970 374294
rect 431206 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 461690 374294
rect 461926 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 492410 374294
rect 492646 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 26490 370894
rect 26726 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 57210 370894
rect 57446 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 87930 370894
rect 88166 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 118650 370894
rect 118886 370658 149370 370894
rect 149606 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 180090 370894
rect 180326 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 210810 370894
rect 211046 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 241530 370894
rect 241766 370658 272250 370894
rect 272486 370658 302970 370894
rect 303206 370658 333690 370894
rect 333926 370658 364410 370894
rect 364646 370658 395130 370894
rect 395366 370658 425850 370894
rect 426086 370658 456570 370894
rect 456806 370658 487290 370894
rect 487526 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 26490 370574
rect 26726 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 57210 370574
rect 57446 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 87930 370574
rect 88166 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 118650 370574
rect 118886 370338 149370 370574
rect 149606 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 180090 370574
rect 180326 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 210810 370574
rect 211046 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 241530 370574
rect 241766 370338 272250 370574
rect 272486 370338 302970 370574
rect 303206 370338 333690 370574
rect 333926 370338 364410 370574
rect 364646 370338 395130 370574
rect 395366 370338 425850 370574
rect 426086 370338 456570 370574
rect 456806 370338 487290 370574
rect 487526 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 21370 367174
rect 21606 366938 52090 367174
rect 52326 366938 82810 367174
rect 83046 366938 113530 367174
rect 113766 366938 144250 367174
rect 144486 366938 174970 367174
rect 175206 366938 205690 367174
rect 205926 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 236410 367174
rect 236646 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 267130 367174
rect 267366 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 297850 367174
rect 298086 366938 328570 367174
rect 328806 366938 359290 367174
rect 359526 366938 390010 367174
rect 390246 366938 420730 367174
rect 420966 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 451450 367174
rect 451686 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 482170 367174
rect 482406 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 21370 366854
rect 21606 366618 52090 366854
rect 52326 366618 82810 366854
rect 83046 366618 113530 366854
rect 113766 366618 144250 366854
rect 144486 366618 174970 366854
rect 175206 366618 205690 366854
rect 205926 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 236410 366854
rect 236646 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 267130 366854
rect 267366 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 297850 366854
rect 298086 366618 328570 366854
rect 328806 366618 359290 366854
rect 359526 366618 390010 366854
rect 390246 366618 420730 366854
rect 420966 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 451450 366854
rect 451686 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 482170 366854
rect 482406 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 16250 363454
rect 16486 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 46970 363454
rect 47206 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 77690 363454
rect 77926 363218 108410 363454
rect 108646 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 139130 363454
rect 139366 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 169850 363454
rect 170086 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 200570 363454
rect 200806 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 231290 363454
rect 231526 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 262010 363454
rect 262246 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 292730 363454
rect 292966 363218 323450 363454
rect 323686 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 354170 363454
rect 354406 363218 384890 363454
rect 385126 363218 415610 363454
rect 415846 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 446330 363454
rect 446566 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 477050 363454
rect 477286 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 507770 363454
rect 508006 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 16250 363134
rect 16486 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 46970 363134
rect 47206 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 77690 363134
rect 77926 362898 108410 363134
rect 108646 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 139130 363134
rect 139366 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 169850 363134
rect 170086 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 200570 363134
rect 200806 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 231290 363134
rect 231526 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 262010 363134
rect 262246 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 292730 363134
rect 292966 362898 323450 363134
rect 323686 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 354170 363134
rect 354406 362898 384890 363134
rect 385126 362898 415610 363134
rect 415846 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 446330 363134
rect 446566 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 477050 363134
rect 477286 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 507770 363134
rect 508006 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 41850 346054
rect 42086 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 72570 346054
rect 72806 345818 103290 346054
rect 103526 345818 134010 346054
rect 134246 345818 164730 346054
rect 164966 345818 195450 346054
rect 195686 345818 226170 346054
rect 226406 345818 256890 346054
rect 257126 345818 287610 346054
rect 287846 345818 318330 346054
rect 318566 345818 349050 346054
rect 349286 345818 379770 346054
rect 380006 345818 410490 346054
rect 410726 345818 441210 346054
rect 441446 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 471930 346054
rect 472166 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 502650 346054
rect 502886 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 41850 345734
rect 42086 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 72570 345734
rect 72806 345498 103290 345734
rect 103526 345498 134010 345734
rect 134246 345498 164730 345734
rect 164966 345498 195450 345734
rect 195686 345498 226170 345734
rect 226406 345498 256890 345734
rect 257126 345498 287610 345734
rect 287846 345498 318330 345734
rect 318566 345498 349050 345734
rect 349286 345498 379770 345734
rect 380006 345498 410490 345734
rect 410726 345498 441210 345734
rect 441446 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 471930 345734
rect 472166 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 502650 345734
rect 502886 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 36730 342334
rect 36966 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 67450 342334
rect 67686 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 98170 342334
rect 98406 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 128890 342334
rect 129126 342098 159610 342334
rect 159846 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 190330 342334
rect 190566 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 221050 342334
rect 221286 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 251770 342334
rect 252006 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 282490 342334
rect 282726 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 313210 342334
rect 313446 342098 343930 342334
rect 344166 342098 374650 342334
rect 374886 342098 405370 342334
rect 405606 342098 436090 342334
rect 436326 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 466810 342334
rect 467046 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 497530 342334
rect 497766 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 36730 342014
rect 36966 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 67450 342014
rect 67686 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 98170 342014
rect 98406 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 128890 342014
rect 129126 341778 159610 342014
rect 159846 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 190330 342014
rect 190566 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 221050 342014
rect 221286 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 251770 342014
rect 252006 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 282490 342014
rect 282726 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 313210 342014
rect 313446 341778 343930 342014
rect 344166 341778 374650 342014
rect 374886 341778 405370 342014
rect 405606 341778 436090 342014
rect 436326 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 466810 342014
rect 467046 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 497530 342014
rect 497766 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 31610 338614
rect 31846 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 62330 338614
rect 62566 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 93050 338614
rect 93286 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 123770 338614
rect 124006 338378 154490 338614
rect 154726 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 185210 338614
rect 185446 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 215930 338614
rect 216166 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 246650 338614
rect 246886 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 277370 338614
rect 277606 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 308090 338614
rect 308326 338378 338810 338614
rect 339046 338378 369530 338614
rect 369766 338378 400250 338614
rect 400486 338378 430970 338614
rect 431206 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 461690 338614
rect 461926 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 492410 338614
rect 492646 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 31610 338294
rect 31846 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 62330 338294
rect 62566 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 93050 338294
rect 93286 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 123770 338294
rect 124006 338058 154490 338294
rect 154726 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 185210 338294
rect 185446 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 215930 338294
rect 216166 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 246650 338294
rect 246886 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 277370 338294
rect 277606 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 308090 338294
rect 308326 338058 338810 338294
rect 339046 338058 369530 338294
rect 369766 338058 400250 338294
rect 400486 338058 430970 338294
rect 431206 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 461690 338294
rect 461926 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 492410 338294
rect 492646 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 26490 334894
rect 26726 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 57210 334894
rect 57446 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 87930 334894
rect 88166 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 118650 334894
rect 118886 334658 149370 334894
rect 149606 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 180090 334894
rect 180326 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 210810 334894
rect 211046 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 241530 334894
rect 241766 334658 272250 334894
rect 272486 334658 302970 334894
rect 303206 334658 333690 334894
rect 333926 334658 364410 334894
rect 364646 334658 395130 334894
rect 395366 334658 425850 334894
rect 426086 334658 456570 334894
rect 456806 334658 487290 334894
rect 487526 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 26490 334574
rect 26726 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 57210 334574
rect 57446 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 87930 334574
rect 88166 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 118650 334574
rect 118886 334338 149370 334574
rect 149606 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 180090 334574
rect 180326 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 210810 334574
rect 211046 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 241530 334574
rect 241766 334338 272250 334574
rect 272486 334338 302970 334574
rect 303206 334338 333690 334574
rect 333926 334338 364410 334574
rect 364646 334338 395130 334574
rect 395366 334338 425850 334574
rect 426086 334338 456570 334574
rect 456806 334338 487290 334574
rect 487526 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 21370 331174
rect 21606 330938 52090 331174
rect 52326 330938 82810 331174
rect 83046 330938 113530 331174
rect 113766 330938 144250 331174
rect 144486 330938 174970 331174
rect 175206 330938 205690 331174
rect 205926 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 236410 331174
rect 236646 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 267130 331174
rect 267366 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 297850 331174
rect 298086 330938 328570 331174
rect 328806 330938 359290 331174
rect 359526 330938 390010 331174
rect 390246 330938 420730 331174
rect 420966 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 451450 331174
rect 451686 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 482170 331174
rect 482406 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 21370 330854
rect 21606 330618 52090 330854
rect 52326 330618 82810 330854
rect 83046 330618 113530 330854
rect 113766 330618 144250 330854
rect 144486 330618 174970 330854
rect 175206 330618 205690 330854
rect 205926 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 236410 330854
rect 236646 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 267130 330854
rect 267366 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 297850 330854
rect 298086 330618 328570 330854
rect 328806 330618 359290 330854
rect 359526 330618 390010 330854
rect 390246 330618 420730 330854
rect 420966 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 451450 330854
rect 451686 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 482170 330854
rect 482406 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 16250 327454
rect 16486 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 46970 327454
rect 47206 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 77690 327454
rect 77926 327218 108410 327454
rect 108646 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 139130 327454
rect 139366 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 169850 327454
rect 170086 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 200570 327454
rect 200806 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 231290 327454
rect 231526 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 262010 327454
rect 262246 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 292730 327454
rect 292966 327218 323450 327454
rect 323686 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 354170 327454
rect 354406 327218 384890 327454
rect 385126 327218 415610 327454
rect 415846 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 446330 327454
rect 446566 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 477050 327454
rect 477286 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 507770 327454
rect 508006 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 16250 327134
rect 16486 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 46970 327134
rect 47206 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 77690 327134
rect 77926 326898 108410 327134
rect 108646 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 139130 327134
rect 139366 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 169850 327134
rect 170086 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 200570 327134
rect 200806 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 231290 327134
rect 231526 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 262010 327134
rect 262246 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 292730 327134
rect 292966 326898 323450 327134
rect 323686 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 354170 327134
rect 354406 326898 384890 327134
rect 385126 326898 415610 327134
rect 415846 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 446330 327134
rect 446566 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 477050 327134
rect 477286 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 507770 327134
rect 508006 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 41850 310054
rect 42086 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 72570 310054
rect 72806 309818 103290 310054
rect 103526 309818 134010 310054
rect 134246 309818 164730 310054
rect 164966 309818 195450 310054
rect 195686 309818 226170 310054
rect 226406 309818 256890 310054
rect 257126 309818 287610 310054
rect 287846 309818 318330 310054
rect 318566 309818 349050 310054
rect 349286 309818 379770 310054
rect 380006 309818 410490 310054
rect 410726 309818 441210 310054
rect 441446 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 471930 310054
rect 472166 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 502650 310054
rect 502886 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 41850 309734
rect 42086 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 72570 309734
rect 72806 309498 103290 309734
rect 103526 309498 134010 309734
rect 134246 309498 164730 309734
rect 164966 309498 195450 309734
rect 195686 309498 226170 309734
rect 226406 309498 256890 309734
rect 257126 309498 287610 309734
rect 287846 309498 318330 309734
rect 318566 309498 349050 309734
rect 349286 309498 379770 309734
rect 380006 309498 410490 309734
rect 410726 309498 441210 309734
rect 441446 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 471930 309734
rect 472166 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 502650 309734
rect 502886 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 36730 306334
rect 36966 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 67450 306334
rect 67686 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 98170 306334
rect 98406 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 128890 306334
rect 129126 306098 159610 306334
rect 159846 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 190330 306334
rect 190566 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 221050 306334
rect 221286 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 251770 306334
rect 252006 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 282490 306334
rect 282726 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 313210 306334
rect 313446 306098 343930 306334
rect 344166 306098 374650 306334
rect 374886 306098 405370 306334
rect 405606 306098 436090 306334
rect 436326 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 466810 306334
rect 467046 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 497530 306334
rect 497766 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 36730 306014
rect 36966 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 67450 306014
rect 67686 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 98170 306014
rect 98406 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 128890 306014
rect 129126 305778 159610 306014
rect 159846 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 190330 306014
rect 190566 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 221050 306014
rect 221286 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 251770 306014
rect 252006 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 282490 306014
rect 282726 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 313210 306014
rect 313446 305778 343930 306014
rect 344166 305778 374650 306014
rect 374886 305778 405370 306014
rect 405606 305778 436090 306014
rect 436326 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 466810 306014
rect 467046 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 497530 306014
rect 497766 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 31610 302614
rect 31846 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 62330 302614
rect 62566 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 93050 302614
rect 93286 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 123770 302614
rect 124006 302378 154490 302614
rect 154726 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 185210 302614
rect 185446 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 215930 302614
rect 216166 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 246650 302614
rect 246886 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 277370 302614
rect 277606 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 308090 302614
rect 308326 302378 338810 302614
rect 339046 302378 369530 302614
rect 369766 302378 400250 302614
rect 400486 302378 430970 302614
rect 431206 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 461690 302614
rect 461926 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 492410 302614
rect 492646 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 31610 302294
rect 31846 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 62330 302294
rect 62566 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 93050 302294
rect 93286 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 123770 302294
rect 124006 302058 154490 302294
rect 154726 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 185210 302294
rect 185446 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 215930 302294
rect 216166 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 246650 302294
rect 246886 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 277370 302294
rect 277606 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 308090 302294
rect 308326 302058 338810 302294
rect 339046 302058 369530 302294
rect 369766 302058 400250 302294
rect 400486 302058 430970 302294
rect 431206 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 461690 302294
rect 461926 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 492410 302294
rect 492646 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 26490 298894
rect 26726 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 57210 298894
rect 57446 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 87930 298894
rect 88166 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 118650 298894
rect 118886 298658 149370 298894
rect 149606 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 180090 298894
rect 180326 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 210810 298894
rect 211046 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 241530 298894
rect 241766 298658 272250 298894
rect 272486 298658 302970 298894
rect 303206 298658 333690 298894
rect 333926 298658 364410 298894
rect 364646 298658 395130 298894
rect 395366 298658 425850 298894
rect 426086 298658 456570 298894
rect 456806 298658 487290 298894
rect 487526 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 26490 298574
rect 26726 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 57210 298574
rect 57446 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 87930 298574
rect 88166 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 118650 298574
rect 118886 298338 149370 298574
rect 149606 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 180090 298574
rect 180326 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 210810 298574
rect 211046 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 241530 298574
rect 241766 298338 272250 298574
rect 272486 298338 302970 298574
rect 303206 298338 333690 298574
rect 333926 298338 364410 298574
rect 364646 298338 395130 298574
rect 395366 298338 425850 298574
rect 426086 298338 456570 298574
rect 456806 298338 487290 298574
rect 487526 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 21370 295174
rect 21606 294938 52090 295174
rect 52326 294938 82810 295174
rect 83046 294938 113530 295174
rect 113766 294938 144250 295174
rect 144486 294938 174970 295174
rect 175206 294938 205690 295174
rect 205926 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 236410 295174
rect 236646 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 267130 295174
rect 267366 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 297850 295174
rect 298086 294938 328570 295174
rect 328806 294938 359290 295174
rect 359526 294938 390010 295174
rect 390246 294938 420730 295174
rect 420966 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 451450 295174
rect 451686 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 482170 295174
rect 482406 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 21370 294854
rect 21606 294618 52090 294854
rect 52326 294618 82810 294854
rect 83046 294618 113530 294854
rect 113766 294618 144250 294854
rect 144486 294618 174970 294854
rect 175206 294618 205690 294854
rect 205926 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 236410 294854
rect 236646 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 267130 294854
rect 267366 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 297850 294854
rect 298086 294618 328570 294854
rect 328806 294618 359290 294854
rect 359526 294618 390010 294854
rect 390246 294618 420730 294854
rect 420966 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 451450 294854
rect 451686 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 482170 294854
rect 482406 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 16250 291454
rect 16486 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 46970 291454
rect 47206 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 77690 291454
rect 77926 291218 108410 291454
rect 108646 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 139130 291454
rect 139366 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 169850 291454
rect 170086 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 200570 291454
rect 200806 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 231290 291454
rect 231526 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 262010 291454
rect 262246 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 292730 291454
rect 292966 291218 323450 291454
rect 323686 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 354170 291454
rect 354406 291218 384890 291454
rect 385126 291218 415610 291454
rect 415846 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 446330 291454
rect 446566 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 477050 291454
rect 477286 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 507770 291454
rect 508006 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 16250 291134
rect 16486 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 46970 291134
rect 47206 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 77690 291134
rect 77926 290898 108410 291134
rect 108646 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 139130 291134
rect 139366 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 169850 291134
rect 170086 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 200570 291134
rect 200806 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 231290 291134
rect 231526 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 262010 291134
rect 262246 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 292730 291134
rect 292966 290898 323450 291134
rect 323686 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 354170 291134
rect 354406 290898 384890 291134
rect 385126 290898 415610 291134
rect 415846 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 446330 291134
rect 446566 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 477050 291134
rect 477286 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 507770 291134
rect 508006 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 276146 277774
rect 276382 277538 276466 277774
rect 276702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 276146 277454
rect 276382 277218 276466 277454
rect 276702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 41850 274054
rect 42086 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 72570 274054
rect 72806 273818 103290 274054
rect 103526 273818 134010 274054
rect 134246 273818 164730 274054
rect 164966 273818 195450 274054
rect 195686 273818 226170 274054
rect 226406 273818 256890 274054
rect 257126 273818 287610 274054
rect 287846 273818 318330 274054
rect 318566 273818 349050 274054
rect 349286 273818 379770 274054
rect 380006 273818 410490 274054
rect 410726 273818 441210 274054
rect 441446 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 471930 274054
rect 472166 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 502650 274054
rect 502886 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 41850 273734
rect 42086 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 72570 273734
rect 72806 273498 103290 273734
rect 103526 273498 134010 273734
rect 134246 273498 164730 273734
rect 164966 273498 195450 273734
rect 195686 273498 226170 273734
rect 226406 273498 256890 273734
rect 257126 273498 287610 273734
rect 287846 273498 318330 273734
rect 318566 273498 349050 273734
rect 349286 273498 379770 273734
rect 380006 273498 410490 273734
rect 410726 273498 441210 273734
rect 441446 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 471930 273734
rect 472166 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 502650 273734
rect 502886 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 36730 270334
rect 36966 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 67450 270334
rect 67686 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 98170 270334
rect 98406 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 128890 270334
rect 129126 270098 159610 270334
rect 159846 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 190330 270334
rect 190566 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 221050 270334
rect 221286 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 251770 270334
rect 252006 270098 268706 270334
rect 268942 270098 269026 270334
rect 269262 270098 282490 270334
rect 282726 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 313210 270334
rect 313446 270098 343930 270334
rect 344166 270098 374650 270334
rect 374886 270098 405370 270334
rect 405606 270098 436090 270334
rect 436326 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 466810 270334
rect 467046 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 497530 270334
rect 497766 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 36730 270014
rect 36966 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 67450 270014
rect 67686 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 98170 270014
rect 98406 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 128890 270014
rect 129126 269778 159610 270014
rect 159846 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 190330 270014
rect 190566 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 221050 270014
rect 221286 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 251770 270014
rect 252006 269778 268706 270014
rect 268942 269778 269026 270014
rect 269262 269778 282490 270014
rect 282726 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 313210 270014
rect 313446 269778 343930 270014
rect 344166 269778 374650 270014
rect 374886 269778 405370 270014
rect 405606 269778 436090 270014
rect 436326 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 466810 270014
rect 467046 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 497530 270014
rect 497766 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 31610 266614
rect 31846 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 62330 266614
rect 62566 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 93050 266614
rect 93286 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 123770 266614
rect 124006 266378 154490 266614
rect 154726 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 185210 266614
rect 185446 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 215930 266614
rect 216166 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 246650 266614
rect 246886 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 277370 266614
rect 277606 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 308090 266614
rect 308326 266378 338810 266614
rect 339046 266378 369530 266614
rect 369766 266378 400250 266614
rect 400486 266378 430970 266614
rect 431206 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 461690 266614
rect 461926 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 492410 266614
rect 492646 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 31610 266294
rect 31846 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 62330 266294
rect 62566 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 93050 266294
rect 93286 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 123770 266294
rect 124006 266058 154490 266294
rect 154726 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 185210 266294
rect 185446 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 215930 266294
rect 216166 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 246650 266294
rect 246886 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 277370 266294
rect 277606 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 308090 266294
rect 308326 266058 338810 266294
rect 339046 266058 369530 266294
rect 369766 266058 400250 266294
rect 400486 266058 430970 266294
rect 431206 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 461690 266294
rect 461926 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 492410 266294
rect 492646 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 26490 262894
rect 26726 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 57210 262894
rect 57446 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 87930 262894
rect 88166 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 118650 262894
rect 118886 262658 149370 262894
rect 149606 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 180090 262894
rect 180326 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 210810 262894
rect 211046 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 241530 262894
rect 241766 262658 272250 262894
rect 272486 262658 302970 262894
rect 303206 262658 333690 262894
rect 333926 262658 364410 262894
rect 364646 262658 395130 262894
rect 395366 262658 425850 262894
rect 426086 262658 456570 262894
rect 456806 262658 487290 262894
rect 487526 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 26490 262574
rect 26726 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 57210 262574
rect 57446 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 87930 262574
rect 88166 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 118650 262574
rect 118886 262338 149370 262574
rect 149606 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 180090 262574
rect 180326 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 210810 262574
rect 211046 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 241530 262574
rect 241766 262338 272250 262574
rect 272486 262338 302970 262574
rect 303206 262338 333690 262574
rect 333926 262338 364410 262574
rect 364646 262338 395130 262574
rect 395366 262338 425850 262574
rect 426086 262338 456570 262574
rect 456806 262338 487290 262574
rect 487526 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 21370 259174
rect 21606 258938 52090 259174
rect 52326 258938 82810 259174
rect 83046 258938 113530 259174
rect 113766 258938 144250 259174
rect 144486 258938 174970 259174
rect 175206 258938 205690 259174
rect 205926 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 236410 259174
rect 236646 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 267130 259174
rect 267366 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 297850 259174
rect 298086 258938 328570 259174
rect 328806 258938 359290 259174
rect 359526 258938 390010 259174
rect 390246 258938 420730 259174
rect 420966 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 451450 259174
rect 451686 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 482170 259174
rect 482406 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 21370 258854
rect 21606 258618 52090 258854
rect 52326 258618 82810 258854
rect 83046 258618 113530 258854
rect 113766 258618 144250 258854
rect 144486 258618 174970 258854
rect 175206 258618 205690 258854
rect 205926 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 236410 258854
rect 236646 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 267130 258854
rect 267366 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 297850 258854
rect 298086 258618 328570 258854
rect 328806 258618 359290 258854
rect 359526 258618 390010 258854
rect 390246 258618 420730 258854
rect 420966 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 451450 258854
rect 451686 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 482170 258854
rect 482406 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 16250 255454
rect 16486 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 46970 255454
rect 47206 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 77690 255454
rect 77926 255218 108410 255454
rect 108646 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 139130 255454
rect 139366 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 169850 255454
rect 170086 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 200570 255454
rect 200806 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 231290 255454
rect 231526 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 262010 255454
rect 262246 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 292730 255454
rect 292966 255218 323450 255454
rect 323686 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 354170 255454
rect 354406 255218 384890 255454
rect 385126 255218 415610 255454
rect 415846 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 446330 255454
rect 446566 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 477050 255454
rect 477286 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 507770 255454
rect 508006 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 16250 255134
rect 16486 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 46970 255134
rect 47206 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 77690 255134
rect 77926 254898 108410 255134
rect 108646 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 139130 255134
rect 139366 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 169850 255134
rect 170086 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 200570 255134
rect 200806 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 231290 255134
rect 231526 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 262010 255134
rect 262246 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 292730 255134
rect 292966 254898 323450 255134
rect 323686 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 354170 255134
rect 354406 254898 384890 255134
rect 385126 254898 415610 255134
rect 415846 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 446330 255134
rect 446566 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 477050 255134
rect 477286 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 507770 255134
rect 508006 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 41850 238054
rect 42086 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 72570 238054
rect 72806 237818 103290 238054
rect 103526 237818 134010 238054
rect 134246 237818 164730 238054
rect 164966 237818 195450 238054
rect 195686 237818 226170 238054
rect 226406 237818 256890 238054
rect 257126 237818 287610 238054
rect 287846 237818 318330 238054
rect 318566 237818 349050 238054
rect 349286 237818 379770 238054
rect 380006 237818 410490 238054
rect 410726 237818 441210 238054
rect 441446 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 471930 238054
rect 472166 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 502650 238054
rect 502886 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 41850 237734
rect 42086 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 72570 237734
rect 72806 237498 103290 237734
rect 103526 237498 134010 237734
rect 134246 237498 164730 237734
rect 164966 237498 195450 237734
rect 195686 237498 226170 237734
rect 226406 237498 256890 237734
rect 257126 237498 287610 237734
rect 287846 237498 318330 237734
rect 318566 237498 349050 237734
rect 349286 237498 379770 237734
rect 380006 237498 410490 237734
rect 410726 237498 441210 237734
rect 441446 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 471930 237734
rect 472166 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 502650 237734
rect 502886 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 36730 234334
rect 36966 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 67450 234334
rect 67686 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 98170 234334
rect 98406 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 128890 234334
rect 129126 234098 159610 234334
rect 159846 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 190330 234334
rect 190566 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 221050 234334
rect 221286 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 251770 234334
rect 252006 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 282490 234334
rect 282726 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 313210 234334
rect 313446 234098 343930 234334
rect 344166 234098 374650 234334
rect 374886 234098 405370 234334
rect 405606 234098 436090 234334
rect 436326 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 466810 234334
rect 467046 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 497530 234334
rect 497766 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 36730 234014
rect 36966 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 67450 234014
rect 67686 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 98170 234014
rect 98406 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 128890 234014
rect 129126 233778 159610 234014
rect 159846 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 190330 234014
rect 190566 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 221050 234014
rect 221286 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 251770 234014
rect 252006 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 282490 234014
rect 282726 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 313210 234014
rect 313446 233778 343930 234014
rect 344166 233778 374650 234014
rect 374886 233778 405370 234014
rect 405606 233778 436090 234014
rect 436326 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 466810 234014
rect 467046 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 497530 234014
rect 497766 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 31610 230614
rect 31846 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 62330 230614
rect 62566 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 93050 230614
rect 93286 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 123770 230614
rect 124006 230378 154490 230614
rect 154726 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 185210 230614
rect 185446 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 215930 230614
rect 216166 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 246650 230614
rect 246886 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 277370 230614
rect 277606 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 308090 230614
rect 308326 230378 338810 230614
rect 339046 230378 369530 230614
rect 369766 230378 400250 230614
rect 400486 230378 430970 230614
rect 431206 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 461690 230614
rect 461926 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 492410 230614
rect 492646 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 31610 230294
rect 31846 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 62330 230294
rect 62566 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 93050 230294
rect 93286 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 123770 230294
rect 124006 230058 154490 230294
rect 154726 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 185210 230294
rect 185446 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 215930 230294
rect 216166 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 246650 230294
rect 246886 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 277370 230294
rect 277606 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 308090 230294
rect 308326 230058 338810 230294
rect 339046 230058 369530 230294
rect 369766 230058 400250 230294
rect 400486 230058 430970 230294
rect 431206 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 461690 230294
rect 461926 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 492410 230294
rect 492646 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 26490 226894
rect 26726 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 57210 226894
rect 57446 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 87930 226894
rect 88166 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 118650 226894
rect 118886 226658 149370 226894
rect 149606 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 180090 226894
rect 180326 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 210810 226894
rect 211046 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 241530 226894
rect 241766 226658 272250 226894
rect 272486 226658 302970 226894
rect 303206 226658 333690 226894
rect 333926 226658 364410 226894
rect 364646 226658 395130 226894
rect 395366 226658 425850 226894
rect 426086 226658 456570 226894
rect 456806 226658 487290 226894
rect 487526 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 26490 226574
rect 26726 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 57210 226574
rect 57446 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 87930 226574
rect 88166 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 118650 226574
rect 118886 226338 149370 226574
rect 149606 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 180090 226574
rect 180326 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 210810 226574
rect 211046 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 241530 226574
rect 241766 226338 272250 226574
rect 272486 226338 302970 226574
rect 303206 226338 333690 226574
rect 333926 226338 364410 226574
rect 364646 226338 395130 226574
rect 395366 226338 425850 226574
rect 426086 226338 456570 226574
rect 456806 226338 487290 226574
rect 487526 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 21370 223174
rect 21606 222938 52090 223174
rect 52326 222938 82810 223174
rect 83046 222938 113530 223174
rect 113766 222938 144250 223174
rect 144486 222938 174970 223174
rect 175206 222938 205690 223174
rect 205926 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 236410 223174
rect 236646 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 267130 223174
rect 267366 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 297850 223174
rect 298086 222938 328570 223174
rect 328806 222938 359290 223174
rect 359526 222938 390010 223174
rect 390246 222938 420730 223174
rect 420966 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 451450 223174
rect 451686 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 482170 223174
rect 482406 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 21370 222854
rect 21606 222618 52090 222854
rect 52326 222618 82810 222854
rect 83046 222618 113530 222854
rect 113766 222618 144250 222854
rect 144486 222618 174970 222854
rect 175206 222618 205690 222854
rect 205926 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 236410 222854
rect 236646 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 267130 222854
rect 267366 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 297850 222854
rect 298086 222618 328570 222854
rect 328806 222618 359290 222854
rect 359526 222618 390010 222854
rect 390246 222618 420730 222854
rect 420966 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 451450 222854
rect 451686 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 482170 222854
rect 482406 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 16250 219454
rect 16486 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 46970 219454
rect 47206 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 77690 219454
rect 77926 219218 108410 219454
rect 108646 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 139130 219454
rect 139366 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 169850 219454
rect 170086 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 200570 219454
rect 200806 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 231290 219454
rect 231526 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 262010 219454
rect 262246 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 292730 219454
rect 292966 219218 323450 219454
rect 323686 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 354170 219454
rect 354406 219218 384890 219454
rect 385126 219218 415610 219454
rect 415846 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 446330 219454
rect 446566 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 477050 219454
rect 477286 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 507770 219454
rect 508006 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 16250 219134
rect 16486 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 46970 219134
rect 47206 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 77690 219134
rect 77926 218898 108410 219134
rect 108646 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 139130 219134
rect 139366 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 169850 219134
rect 170086 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 200570 219134
rect 200806 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 231290 219134
rect 231526 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 262010 219134
rect 262246 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 292730 219134
rect 292966 218898 323450 219134
rect 323686 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 354170 219134
rect 354406 218898 384890 219134
rect 385126 218898 415610 219134
rect 415846 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 446330 219134
rect 446566 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 477050 219134
rect 477286 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 507770 219134
rect 508006 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 41850 202054
rect 42086 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 72570 202054
rect 72806 201818 103290 202054
rect 103526 201818 134010 202054
rect 134246 201818 164730 202054
rect 164966 201818 195450 202054
rect 195686 201818 226170 202054
rect 226406 201818 256890 202054
rect 257126 201818 287610 202054
rect 287846 201818 318330 202054
rect 318566 201818 349050 202054
rect 349286 201818 379770 202054
rect 380006 201818 410490 202054
rect 410726 201818 441210 202054
rect 441446 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 471930 202054
rect 472166 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 502650 202054
rect 502886 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 41850 201734
rect 42086 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 72570 201734
rect 72806 201498 103290 201734
rect 103526 201498 134010 201734
rect 134246 201498 164730 201734
rect 164966 201498 195450 201734
rect 195686 201498 226170 201734
rect 226406 201498 256890 201734
rect 257126 201498 287610 201734
rect 287846 201498 318330 201734
rect 318566 201498 349050 201734
rect 349286 201498 379770 201734
rect 380006 201498 410490 201734
rect 410726 201498 441210 201734
rect 441446 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 471930 201734
rect 472166 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 502650 201734
rect 502886 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 36730 198334
rect 36966 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 67450 198334
rect 67686 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 98170 198334
rect 98406 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 128890 198334
rect 129126 198098 159610 198334
rect 159846 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 190330 198334
rect 190566 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 221050 198334
rect 221286 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 251770 198334
rect 252006 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 282490 198334
rect 282726 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 313210 198334
rect 313446 198098 343930 198334
rect 344166 198098 374650 198334
rect 374886 198098 436090 198334
rect 436326 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 466810 198334
rect 467046 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 497530 198334
rect 497766 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 36730 198014
rect 36966 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 67450 198014
rect 67686 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 98170 198014
rect 98406 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 128890 198014
rect 129126 197778 159610 198014
rect 159846 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 190330 198014
rect 190566 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 221050 198014
rect 221286 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 251770 198014
rect 252006 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 282490 198014
rect 282726 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 313210 198014
rect 313446 197778 343930 198014
rect 344166 197778 374650 198014
rect 374886 197778 436090 198014
rect 436326 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 466810 198014
rect 467046 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 497530 198014
rect 497766 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 31610 194614
rect 31846 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 62330 194614
rect 62566 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 93050 194614
rect 93286 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 123770 194614
rect 124006 194378 154490 194614
rect 154726 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 185210 194614
rect 185446 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 215930 194614
rect 216166 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 246650 194614
rect 246886 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 277370 194614
rect 277606 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 308090 194614
rect 308326 194378 338810 194614
rect 339046 194378 369530 194614
rect 369766 194431 430970 194614
rect 369766 194378 400250 194431
rect -8726 194294 400250 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 31610 194294
rect 31846 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 62330 194294
rect 62566 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 93050 194294
rect 93286 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 123770 194294
rect 124006 194058 154490 194294
rect 154726 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 185210 194294
rect 185446 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 215930 194294
rect 216166 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 246650 194294
rect 246886 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 277370 194294
rect 277606 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 308090 194294
rect 308326 194058 338810 194294
rect 339046 194058 369530 194294
rect 369766 194195 400250 194294
rect 400486 194378 430970 194431
rect 431206 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 461690 194614
rect 461926 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 492410 194614
rect 492646 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect 400486 194294 592650 194378
rect 400486 194195 430970 194294
rect 369766 194058 430970 194195
rect 431206 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 461690 194294
rect 461926 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 492410 194294
rect 492646 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 26490 190894
rect 26726 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 57210 190894
rect 57446 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 87930 190894
rect 88166 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 118650 190894
rect 118886 190658 149370 190894
rect 149606 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 180090 190894
rect 180326 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 210810 190894
rect 211046 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 241530 190894
rect 241766 190658 272250 190894
rect 272486 190658 302970 190894
rect 303206 190658 333690 190894
rect 333926 190658 364410 190894
rect 364646 190658 395130 190894
rect 395366 190658 425850 190894
rect 426086 190658 456570 190894
rect 456806 190658 487290 190894
rect 487526 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 26490 190574
rect 26726 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 57210 190574
rect 57446 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 87930 190574
rect 88166 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 118650 190574
rect 118886 190338 149370 190574
rect 149606 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 180090 190574
rect 180326 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 210810 190574
rect 211046 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 241530 190574
rect 241766 190338 272250 190574
rect 272486 190338 302970 190574
rect 303206 190338 333690 190574
rect 333926 190338 364410 190574
rect 364646 190338 395130 190574
rect 395366 190338 425850 190574
rect 426086 190338 456570 190574
rect 456806 190338 487290 190574
rect 487526 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 21370 187174
rect 21606 186938 52090 187174
rect 52326 186938 82810 187174
rect 83046 186938 113530 187174
rect 113766 186938 144250 187174
rect 144486 186938 174970 187174
rect 175206 186938 205690 187174
rect 205926 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 236410 187174
rect 236646 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 267130 187174
rect 267366 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 297850 187174
rect 298086 186938 328570 187174
rect 328806 186938 359290 187174
rect 359526 186938 390010 187174
rect 390246 186938 420730 187174
rect 420966 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 451450 187174
rect 451686 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 482170 187174
rect 482406 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 21370 186854
rect 21606 186618 52090 186854
rect 52326 186618 82810 186854
rect 83046 186618 113530 186854
rect 113766 186618 144250 186854
rect 144486 186618 174970 186854
rect 175206 186618 205690 186854
rect 205926 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 236410 186854
rect 236646 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 267130 186854
rect 267366 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 297850 186854
rect 298086 186618 328570 186854
rect 328806 186618 359290 186854
rect 359526 186618 390010 186854
rect 390246 186618 420730 186854
rect 420966 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 451450 186854
rect 451686 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 482170 186854
rect 482406 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 16250 183454
rect 16486 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 46970 183454
rect 47206 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 139130 183454
rect 139366 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 169850 183454
rect 170086 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 200570 183454
rect 200806 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 231290 183454
rect 231526 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 262010 183454
rect 262246 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 292730 183454
rect 292966 183218 323450 183454
rect 323686 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 354170 183454
rect 354406 183218 384890 183454
rect 385126 183218 415610 183454
rect 415846 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 446330 183454
rect 446566 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 477050 183454
rect 477286 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 507770 183454
rect 508006 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 16250 183134
rect 16486 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 46970 183134
rect 47206 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 139130 183134
rect 139366 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 169850 183134
rect 170086 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 200570 183134
rect 200806 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 231290 183134
rect 231526 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 262010 183134
rect 262246 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 292730 183134
rect 292966 182898 323450 183134
rect 323686 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 354170 183134
rect 354406 182898 384890 183134
rect 385126 182898 415610 183134
rect 415846 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 446330 183134
rect 446566 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 477050 183134
rect 477286 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 507770 183134
rect 508006 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 41850 166054
rect 42086 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 72570 166054
rect 72806 165818 103290 166054
rect 103526 165818 134010 166054
rect 134246 165818 164730 166054
rect 164966 165818 195450 166054
rect 195686 165818 226170 166054
rect 226406 165818 256890 166054
rect 257126 165818 287610 166054
rect 287846 165818 318330 166054
rect 318566 165818 349050 166054
rect 349286 165818 379770 166054
rect 380006 165818 410490 166054
rect 410726 165818 441210 166054
rect 441446 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 471930 166054
rect 472166 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 502650 166054
rect 502886 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 41850 165734
rect 42086 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 72570 165734
rect 72806 165498 103290 165734
rect 103526 165498 134010 165734
rect 134246 165498 164730 165734
rect 164966 165498 195450 165734
rect 195686 165498 226170 165734
rect 226406 165498 256890 165734
rect 257126 165498 287610 165734
rect 287846 165498 318330 165734
rect 318566 165498 349050 165734
rect 349286 165498 379770 165734
rect 380006 165498 410490 165734
rect 410726 165498 441210 165734
rect 441446 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 471930 165734
rect 472166 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 502650 165734
rect 502886 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 36730 162334
rect 36966 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 67450 162334
rect 67686 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 98170 162334
rect 98406 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 128890 162334
rect 129126 162098 159610 162334
rect 159846 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 190330 162334
rect 190566 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 221050 162334
rect 221286 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 251770 162334
rect 252006 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 282490 162334
rect 282726 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 313210 162334
rect 313446 162098 343930 162334
rect 344166 162098 374650 162334
rect 374886 162098 405370 162334
rect 405606 162098 436090 162334
rect 436326 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 466810 162334
rect 467046 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 497530 162334
rect 497766 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 36730 162014
rect 36966 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 67450 162014
rect 67686 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 98170 162014
rect 98406 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 128890 162014
rect 129126 161778 159610 162014
rect 159846 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 190330 162014
rect 190566 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 221050 162014
rect 221286 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 251770 162014
rect 252006 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 282490 162014
rect 282726 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 313210 162014
rect 313446 161778 343930 162014
rect 344166 161778 374650 162014
rect 374886 161778 405370 162014
rect 405606 161778 436090 162014
rect 436326 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 466810 162014
rect 467046 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 497530 162014
rect 497766 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 31610 158614
rect 31846 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 62330 158614
rect 62566 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 93050 158614
rect 93286 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 123770 158614
rect 124006 158378 154490 158614
rect 154726 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 185210 158614
rect 185446 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 215930 158614
rect 216166 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 246650 158614
rect 246886 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 277370 158614
rect 277606 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 308090 158614
rect 308326 158378 338810 158614
rect 339046 158378 369530 158614
rect 369766 158378 400250 158614
rect 400486 158378 430970 158614
rect 431206 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 461690 158614
rect 461926 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 492410 158614
rect 492646 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 31610 158294
rect 31846 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 62330 158294
rect 62566 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 93050 158294
rect 93286 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 123770 158294
rect 124006 158058 154490 158294
rect 154726 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 185210 158294
rect 185446 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 215930 158294
rect 216166 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 246650 158294
rect 246886 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 277370 158294
rect 277606 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 308090 158294
rect 308326 158058 338810 158294
rect 339046 158058 369530 158294
rect 369766 158058 400250 158294
rect 400486 158058 430970 158294
rect 431206 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 461690 158294
rect 461926 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 492410 158294
rect 492646 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 26490 154894
rect 26726 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 57210 154894
rect 57446 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 87930 154894
rect 88166 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 118650 154894
rect 118886 154658 149370 154894
rect 149606 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 180090 154894
rect 180326 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 210810 154894
rect 211046 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 241530 154894
rect 241766 154658 272250 154894
rect 272486 154658 302970 154894
rect 303206 154658 333690 154894
rect 333926 154658 364410 154894
rect 364646 154658 395130 154894
rect 395366 154658 425850 154894
rect 426086 154658 456570 154894
rect 456806 154658 487290 154894
rect 487526 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 26490 154574
rect 26726 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 57210 154574
rect 57446 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 87930 154574
rect 88166 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 118650 154574
rect 118886 154338 149370 154574
rect 149606 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 180090 154574
rect 180326 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 210810 154574
rect 211046 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 241530 154574
rect 241766 154338 272250 154574
rect 272486 154338 302970 154574
rect 303206 154338 333690 154574
rect 333926 154338 364410 154574
rect 364646 154338 395130 154574
rect 395366 154338 425850 154574
rect 426086 154338 456570 154574
rect 456806 154338 487290 154574
rect 487526 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 21370 151174
rect 21606 150938 52090 151174
rect 52326 150938 82810 151174
rect 83046 150938 113530 151174
rect 113766 150938 144250 151174
rect 144486 150938 174970 151174
rect 175206 150938 205690 151174
rect 205926 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 236410 151174
rect 236646 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 267130 151174
rect 267366 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 297850 151174
rect 298086 150938 328570 151174
rect 328806 150938 359290 151174
rect 359526 150938 390010 151174
rect 390246 150938 420730 151174
rect 420966 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 451450 151174
rect 451686 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 482170 151174
rect 482406 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 21370 150854
rect 21606 150618 52090 150854
rect 52326 150618 82810 150854
rect 83046 150618 113530 150854
rect 113766 150618 144250 150854
rect 144486 150618 174970 150854
rect 175206 150618 205690 150854
rect 205926 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 236410 150854
rect 236646 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 267130 150854
rect 267366 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 297850 150854
rect 298086 150618 328570 150854
rect 328806 150618 359290 150854
rect 359526 150618 390010 150854
rect 390246 150618 420730 150854
rect 420966 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 451450 150854
rect 451686 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 482170 150854
rect 482406 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 16250 147454
rect 16486 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 46970 147454
rect 47206 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 139130 147454
rect 139366 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 169850 147454
rect 170086 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 200570 147454
rect 200806 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 231290 147454
rect 231526 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 262010 147454
rect 262246 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 292730 147454
rect 292966 147218 323450 147454
rect 323686 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 354170 147454
rect 354406 147218 384890 147454
rect 385126 147218 415610 147454
rect 415846 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 446330 147454
rect 446566 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 477050 147454
rect 477286 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 507770 147454
rect 508006 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 16250 147134
rect 16486 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 46970 147134
rect 47206 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 139130 147134
rect 139366 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 169850 147134
rect 170086 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 200570 147134
rect 200806 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 231290 147134
rect 231526 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 262010 147134
rect 262246 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 292730 147134
rect 292966 146898 323450 147134
rect 323686 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 354170 147134
rect 354406 146898 384890 147134
rect 385126 146898 415610 147134
rect 415846 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 446330 147134
rect 446566 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 477050 147134
rect 477286 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 507770 147134
rect 508006 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 41850 130054
rect 42086 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 72570 130054
rect 72806 129818 103290 130054
rect 103526 129818 134010 130054
rect 134246 129818 164730 130054
rect 164966 129818 195450 130054
rect 195686 129818 226170 130054
rect 226406 129818 256890 130054
rect 257126 129818 287610 130054
rect 287846 129818 318330 130054
rect 318566 129818 349050 130054
rect 349286 129818 379770 130054
rect 380006 129818 410490 130054
rect 410726 129818 441210 130054
rect 441446 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 471930 130054
rect 472166 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 502650 130054
rect 502886 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 41850 129734
rect 42086 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 72570 129734
rect 72806 129498 103290 129734
rect 103526 129498 134010 129734
rect 134246 129498 164730 129734
rect 164966 129498 195450 129734
rect 195686 129498 226170 129734
rect 226406 129498 256890 129734
rect 257126 129498 287610 129734
rect 287846 129498 318330 129734
rect 318566 129498 349050 129734
rect 349286 129498 379770 129734
rect 380006 129498 410490 129734
rect 410726 129498 441210 129734
rect 441446 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 471930 129734
rect 472166 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 502650 129734
rect 502886 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 36730 126334
rect 36966 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 67450 126334
rect 67686 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 98170 126334
rect 98406 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 128890 126334
rect 129126 126098 159610 126334
rect 159846 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 190330 126334
rect 190566 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 221050 126334
rect 221286 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 251770 126334
rect 252006 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 282490 126334
rect 282726 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 313210 126334
rect 313446 126098 343930 126334
rect 344166 126098 374650 126334
rect 374886 126098 405370 126334
rect 405606 126098 436090 126334
rect 436326 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 466810 126334
rect 467046 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 497530 126334
rect 497766 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 36730 126014
rect 36966 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 67450 126014
rect 67686 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 98170 126014
rect 98406 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 128890 126014
rect 129126 125778 159610 126014
rect 159846 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 190330 126014
rect 190566 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 221050 126014
rect 221286 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 251770 126014
rect 252006 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 282490 126014
rect 282726 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 313210 126014
rect 313446 125778 343930 126014
rect 344166 125778 374650 126014
rect 374886 125778 405370 126014
rect 405606 125778 436090 126014
rect 436326 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 466810 126014
rect 467046 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 497530 126014
rect 497766 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 31610 122614
rect 31846 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 62330 122614
rect 62566 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 93050 122614
rect 93286 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 123770 122614
rect 124006 122378 154490 122614
rect 154726 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 185210 122614
rect 185446 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 215930 122614
rect 216166 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 246650 122614
rect 246886 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 277370 122614
rect 277606 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 308090 122614
rect 308326 122378 338810 122614
rect 339046 122378 369530 122614
rect 369766 122378 400250 122614
rect 400486 122378 430970 122614
rect 431206 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 461690 122614
rect 461926 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 492410 122614
rect 492646 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 31610 122294
rect 31846 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 62330 122294
rect 62566 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 93050 122294
rect 93286 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 123770 122294
rect 124006 122058 154490 122294
rect 154726 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 185210 122294
rect 185446 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 215930 122294
rect 216166 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 246650 122294
rect 246886 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 277370 122294
rect 277606 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 308090 122294
rect 308326 122058 338810 122294
rect 339046 122058 369530 122294
rect 369766 122058 400250 122294
rect 400486 122058 430970 122294
rect 431206 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 461690 122294
rect 461926 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 492410 122294
rect 492646 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 26490 118894
rect 26726 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 57210 118894
rect 57446 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 87930 118894
rect 88166 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 118650 118894
rect 118886 118658 149370 118894
rect 149606 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 180090 118894
rect 180326 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 210810 118894
rect 211046 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 241530 118894
rect 241766 118658 272250 118894
rect 272486 118658 302970 118894
rect 303206 118658 333690 118894
rect 333926 118658 364410 118894
rect 364646 118658 395130 118894
rect 395366 118658 425850 118894
rect 426086 118658 456570 118894
rect 456806 118658 487290 118894
rect 487526 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 26490 118574
rect 26726 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 57210 118574
rect 57446 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 87930 118574
rect 88166 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 118650 118574
rect 118886 118338 149370 118574
rect 149606 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 180090 118574
rect 180326 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 210810 118574
rect 211046 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 241530 118574
rect 241766 118338 272250 118574
rect 272486 118338 302970 118574
rect 303206 118338 333690 118574
rect 333926 118338 364410 118574
rect 364646 118338 395130 118574
rect 395366 118338 425850 118574
rect 426086 118338 456570 118574
rect 456806 118338 487290 118574
rect 487526 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 21370 115174
rect 21606 114938 52090 115174
rect 52326 114938 82810 115174
rect 83046 114938 113530 115174
rect 113766 114938 144250 115174
rect 144486 114938 174970 115174
rect 175206 114938 205690 115174
rect 205926 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 236410 115174
rect 236646 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 267130 115174
rect 267366 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 297850 115174
rect 298086 114938 328570 115174
rect 328806 114938 359290 115174
rect 359526 114938 390010 115174
rect 390246 114938 420730 115174
rect 420966 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 451450 115174
rect 451686 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 482170 115174
rect 482406 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 21370 114854
rect 21606 114618 52090 114854
rect 52326 114618 82810 114854
rect 83046 114618 113530 114854
rect 113766 114618 144250 114854
rect 144486 114618 174970 114854
rect 175206 114618 205690 114854
rect 205926 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 236410 114854
rect 236646 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 267130 114854
rect 267366 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 297850 114854
rect 298086 114618 328570 114854
rect 328806 114618 359290 114854
rect 359526 114618 390010 114854
rect 390246 114618 420730 114854
rect 420966 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 451450 114854
rect 451686 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 482170 114854
rect 482406 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 16250 111454
rect 16486 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 46970 111454
rect 47206 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 139130 111454
rect 139366 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 169850 111454
rect 170086 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 200570 111454
rect 200806 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 231290 111454
rect 231526 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 262010 111454
rect 262246 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 292730 111454
rect 292966 111218 323450 111454
rect 323686 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 354170 111454
rect 354406 111218 384890 111454
rect 385126 111218 415610 111454
rect 415846 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 446330 111454
rect 446566 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 477050 111454
rect 477286 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 507770 111454
rect 508006 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 16250 111134
rect 16486 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 46970 111134
rect 47206 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 139130 111134
rect 139366 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 169850 111134
rect 170086 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 200570 111134
rect 200806 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 231290 111134
rect 231526 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 262010 111134
rect 262246 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 292730 111134
rect 292966 110898 323450 111134
rect 323686 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 354170 111134
rect 354406 110898 384890 111134
rect 385126 110898 415610 111134
rect 415846 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 446330 111134
rect 446566 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 477050 111134
rect 477286 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 507770 111134
rect 508006 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 41850 94054
rect 42086 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 72570 94054
rect 72806 93818 103290 94054
rect 103526 93818 134010 94054
rect 134246 93818 164730 94054
rect 164966 93818 195450 94054
rect 195686 93818 226170 94054
rect 226406 93818 256890 94054
rect 257126 93818 287610 94054
rect 287846 93818 318330 94054
rect 318566 93818 349050 94054
rect 349286 93818 379770 94054
rect 380006 93818 410490 94054
rect 410726 93818 441210 94054
rect 441446 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 471930 94054
rect 472166 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 502650 94054
rect 502886 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 41850 93734
rect 42086 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 72570 93734
rect 72806 93498 103290 93734
rect 103526 93498 134010 93734
rect 134246 93498 164730 93734
rect 164966 93498 195450 93734
rect 195686 93498 226170 93734
rect 226406 93498 256890 93734
rect 257126 93498 287610 93734
rect 287846 93498 318330 93734
rect 318566 93498 349050 93734
rect 349286 93498 379770 93734
rect 380006 93498 410490 93734
rect 410726 93498 441210 93734
rect 441446 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 471930 93734
rect 472166 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 502650 93734
rect 502886 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 36730 90334
rect 36966 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 67450 90334
rect 67686 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 98170 90334
rect 98406 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 128890 90334
rect 129126 90098 159610 90334
rect 159846 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 190330 90334
rect 190566 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 221050 90334
rect 221286 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 251770 90334
rect 252006 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 282490 90334
rect 282726 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 313210 90334
rect 313446 90098 343930 90334
rect 344166 90098 374650 90334
rect 374886 90098 405370 90334
rect 405606 90098 436090 90334
rect 436326 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 466810 90334
rect 467046 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 497530 90334
rect 497766 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 36730 90014
rect 36966 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 67450 90014
rect 67686 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 98170 90014
rect 98406 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 128890 90014
rect 129126 89778 159610 90014
rect 159846 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 190330 90014
rect 190566 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 221050 90014
rect 221286 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 251770 90014
rect 252006 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 282490 90014
rect 282726 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 313210 90014
rect 313446 89778 343930 90014
rect 344166 89778 374650 90014
rect 374886 89778 405370 90014
rect 405606 89778 436090 90014
rect 436326 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 466810 90014
rect 467046 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 497530 90014
rect 497766 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 31610 86614
rect 31846 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 62330 86614
rect 62566 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 93050 86614
rect 93286 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 123770 86614
rect 124006 86378 154490 86614
rect 154726 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 185210 86614
rect 185446 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 215930 86614
rect 216166 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 246650 86614
rect 246886 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 277370 86614
rect 277606 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 308090 86614
rect 308326 86378 338810 86614
rect 339046 86378 369530 86614
rect 369766 86378 400250 86614
rect 400486 86378 430970 86614
rect 431206 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 461690 86614
rect 461926 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 492410 86614
rect 492646 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 31610 86294
rect 31846 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 62330 86294
rect 62566 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 93050 86294
rect 93286 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 123770 86294
rect 124006 86058 154490 86294
rect 154726 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 185210 86294
rect 185446 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 215930 86294
rect 216166 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 246650 86294
rect 246886 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 277370 86294
rect 277606 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 308090 86294
rect 308326 86058 338810 86294
rect 339046 86058 369530 86294
rect 369766 86058 400250 86294
rect 400486 86058 430970 86294
rect 431206 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 461690 86294
rect 461926 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 492410 86294
rect 492646 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 26490 82894
rect 26726 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 57210 82894
rect 57446 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 87930 82894
rect 88166 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 118650 82894
rect 118886 82658 149370 82894
rect 149606 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 180090 82894
rect 180326 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 210810 82894
rect 211046 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 241530 82894
rect 241766 82658 272250 82894
rect 272486 82658 302970 82894
rect 303206 82658 333690 82894
rect 333926 82658 364410 82894
rect 364646 82658 395130 82894
rect 395366 82658 425850 82894
rect 426086 82658 456570 82894
rect 456806 82658 487290 82894
rect 487526 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 26490 82574
rect 26726 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 57210 82574
rect 57446 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 87930 82574
rect 88166 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 118650 82574
rect 118886 82338 149370 82574
rect 149606 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 180090 82574
rect 180326 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 210810 82574
rect 211046 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 241530 82574
rect 241766 82338 272250 82574
rect 272486 82338 302970 82574
rect 303206 82338 333690 82574
rect 333926 82338 364410 82574
rect 364646 82338 395130 82574
rect 395366 82338 425850 82574
rect 426086 82338 456570 82574
rect 456806 82338 487290 82574
rect 487526 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 21370 79174
rect 21606 78938 52090 79174
rect 52326 78938 82810 79174
rect 83046 78938 113530 79174
rect 113766 78938 144250 79174
rect 144486 78938 174970 79174
rect 175206 78938 205690 79174
rect 205926 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 236410 79174
rect 236646 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 267130 79174
rect 267366 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 297850 79174
rect 298086 78938 328570 79174
rect 328806 78938 359290 79174
rect 359526 78938 390010 79174
rect 390246 78938 420730 79174
rect 420966 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 451450 79174
rect 451686 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 482170 79174
rect 482406 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 21370 78854
rect 21606 78618 52090 78854
rect 52326 78618 82810 78854
rect 83046 78618 113530 78854
rect 113766 78618 144250 78854
rect 144486 78618 174970 78854
rect 175206 78618 205690 78854
rect 205926 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 236410 78854
rect 236646 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 267130 78854
rect 267366 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 297850 78854
rect 298086 78618 328570 78854
rect 328806 78618 359290 78854
rect 359526 78618 390010 78854
rect 390246 78618 420730 78854
rect 420966 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 451450 78854
rect 451686 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 482170 78854
rect 482406 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 16250 75454
rect 16486 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 46970 75454
rect 47206 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 139130 75454
rect 139366 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 169850 75454
rect 170086 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 200570 75454
rect 200806 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 231290 75454
rect 231526 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 262010 75454
rect 262246 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 292730 75454
rect 292966 75218 323450 75454
rect 323686 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 354170 75454
rect 354406 75218 384890 75454
rect 385126 75218 415610 75454
rect 415846 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 446330 75454
rect 446566 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 477050 75454
rect 477286 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 507770 75454
rect 508006 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 16250 75134
rect 16486 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 46970 75134
rect 47206 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 139130 75134
rect 139366 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 169850 75134
rect 170086 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 200570 75134
rect 200806 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 231290 75134
rect 231526 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 262010 75134
rect 262246 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 292730 75134
rect 292966 74898 323450 75134
rect 323686 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 354170 75134
rect 354406 74898 384890 75134
rect 385126 74898 415610 75134
rect 415846 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 446330 75134
rect 446566 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 477050 75134
rect 477286 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 507770 75134
rect 508006 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 41850 58054
rect 42086 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 72570 58054
rect 72806 57818 103290 58054
rect 103526 57818 134010 58054
rect 134246 57818 164730 58054
rect 164966 57818 195450 58054
rect 195686 57818 226170 58054
rect 226406 57818 256890 58054
rect 257126 57818 287610 58054
rect 287846 57818 318330 58054
rect 318566 57818 349050 58054
rect 349286 57818 379770 58054
rect 380006 57818 410490 58054
rect 410726 57818 441210 58054
rect 441446 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 471930 58054
rect 472166 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 502650 58054
rect 502886 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 41850 57734
rect 42086 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 72570 57734
rect 72806 57498 103290 57734
rect 103526 57498 134010 57734
rect 134246 57498 164730 57734
rect 164966 57498 195450 57734
rect 195686 57498 226170 57734
rect 226406 57498 256890 57734
rect 257126 57498 287610 57734
rect 287846 57498 318330 57734
rect 318566 57498 349050 57734
rect 349286 57498 379770 57734
rect 380006 57498 410490 57734
rect 410726 57498 441210 57734
rect 441446 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 471930 57734
rect 472166 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 502650 57734
rect 502886 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 36730 54334
rect 36966 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 67450 54334
rect 67686 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 98170 54334
rect 98406 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 128890 54334
rect 129126 54098 159610 54334
rect 159846 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 190330 54334
rect 190566 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 221050 54334
rect 221286 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 251770 54334
rect 252006 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 282490 54334
rect 282726 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 313210 54334
rect 313446 54098 343930 54334
rect 344166 54098 374650 54334
rect 374886 54098 405370 54334
rect 405606 54098 436090 54334
rect 436326 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 466810 54334
rect 467046 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 497530 54334
rect 497766 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 36730 54014
rect 36966 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 67450 54014
rect 67686 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 98170 54014
rect 98406 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 128890 54014
rect 129126 53778 159610 54014
rect 159846 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 190330 54014
rect 190566 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 221050 54014
rect 221286 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 251770 54014
rect 252006 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 282490 54014
rect 282726 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 313210 54014
rect 313446 53778 343930 54014
rect 344166 53778 374650 54014
rect 374886 53778 405370 54014
rect 405606 53778 436090 54014
rect 436326 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 466810 54014
rect 467046 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 497530 54014
rect 497766 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 31610 50614
rect 31846 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 62330 50614
rect 62566 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 93050 50614
rect 93286 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 123770 50614
rect 124006 50378 154490 50614
rect 154726 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 185210 50614
rect 185446 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 215930 50614
rect 216166 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 246650 50614
rect 246886 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 277370 50614
rect 277606 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 308090 50614
rect 308326 50378 338810 50614
rect 339046 50378 369530 50614
rect 369766 50378 400250 50614
rect 400486 50378 430970 50614
rect 431206 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 461690 50614
rect 461926 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 492410 50614
rect 492646 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 31610 50294
rect 31846 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 62330 50294
rect 62566 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 93050 50294
rect 93286 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 123770 50294
rect 124006 50058 154490 50294
rect 154726 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 185210 50294
rect 185446 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 215930 50294
rect 216166 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 246650 50294
rect 246886 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 277370 50294
rect 277606 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 308090 50294
rect 308326 50058 338810 50294
rect 339046 50058 369530 50294
rect 369766 50058 400250 50294
rect 400486 50058 430970 50294
rect 431206 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 461690 50294
rect 461926 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 492410 50294
rect 492646 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 26490 46894
rect 26726 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 57210 46894
rect 57446 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 87930 46894
rect 88166 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 118650 46894
rect 118886 46658 149370 46894
rect 149606 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 180090 46894
rect 180326 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 210810 46894
rect 211046 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 241530 46894
rect 241766 46658 272250 46894
rect 272486 46658 302970 46894
rect 303206 46658 333690 46894
rect 333926 46658 364410 46894
rect 364646 46658 395130 46894
rect 395366 46658 425850 46894
rect 426086 46658 456570 46894
rect 456806 46658 487290 46894
rect 487526 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 26490 46574
rect 26726 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 57210 46574
rect 57446 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 87930 46574
rect 88166 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 118650 46574
rect 118886 46338 149370 46574
rect 149606 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 180090 46574
rect 180326 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 210810 46574
rect 211046 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 241530 46574
rect 241766 46338 272250 46574
rect 272486 46338 302970 46574
rect 303206 46338 333690 46574
rect 333926 46338 364410 46574
rect 364646 46338 395130 46574
rect 395366 46338 425850 46574
rect 426086 46338 456570 46574
rect 456806 46338 487290 46574
rect 487526 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 21370 43174
rect 21606 42938 52090 43174
rect 52326 42938 82810 43174
rect 83046 42938 113530 43174
rect 113766 42938 144250 43174
rect 144486 42938 174970 43174
rect 175206 42938 205690 43174
rect 205926 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 236410 43174
rect 236646 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 267130 43174
rect 267366 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 297850 43174
rect 298086 42938 328570 43174
rect 328806 42938 359290 43174
rect 359526 42938 390010 43174
rect 390246 42938 420730 43174
rect 420966 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 451450 43174
rect 451686 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 482170 43174
rect 482406 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 21370 42854
rect 21606 42618 52090 42854
rect 52326 42618 82810 42854
rect 83046 42618 113530 42854
rect 113766 42618 144250 42854
rect 144486 42618 174970 42854
rect 175206 42618 205690 42854
rect 205926 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 236410 42854
rect 236646 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 267130 42854
rect 267366 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 297850 42854
rect 298086 42618 328570 42854
rect 328806 42618 359290 42854
rect 359526 42618 390010 42854
rect 390246 42618 420730 42854
rect 420966 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 451450 42854
rect 451686 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 482170 42854
rect 482406 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 16250 39454
rect 16486 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 46970 39454
rect 47206 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 139130 39454
rect 139366 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 169850 39454
rect 170086 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 200570 39454
rect 200806 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 231290 39454
rect 231526 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 262010 39454
rect 262246 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 292730 39454
rect 292966 39218 323450 39454
rect 323686 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 354170 39454
rect 354406 39218 384890 39454
rect 385126 39218 415610 39454
rect 415846 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 446330 39454
rect 446566 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 477050 39454
rect 477286 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 507770 39454
rect 508006 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 16250 39134
rect 16486 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 46970 39134
rect 47206 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 139130 39134
rect 139366 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 169850 39134
rect 170086 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 200570 39134
rect 200806 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 231290 39134
rect 231526 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 262010 39134
rect 262246 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 292730 39134
rect 292966 38898 323450 39134
rect 323686 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 354170 39134
rect 354406 38898 384890 39134
rect 385126 38898 415610 39134
rect 415846 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 446330 39134
rect 446566 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 477050 39134
rect 477286 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 507770 39134
rect 508006 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 41850 22054
rect 42086 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 72570 22054
rect 72806 21818 103290 22054
rect 103526 21818 134010 22054
rect 134246 21818 164730 22054
rect 164966 21818 195450 22054
rect 195686 21818 226170 22054
rect 226406 21818 256890 22054
rect 257126 21818 287610 22054
rect 287846 21818 318330 22054
rect 318566 21818 349050 22054
rect 349286 21818 379770 22054
rect 380006 21818 410490 22054
rect 410726 21818 441210 22054
rect 441446 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 471930 22054
rect 472166 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 502650 22054
rect 502886 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 41850 21734
rect 42086 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 72570 21734
rect 72806 21498 103290 21734
rect 103526 21498 134010 21734
rect 134246 21498 164730 21734
rect 164966 21498 195450 21734
rect 195686 21498 226170 21734
rect 226406 21498 256890 21734
rect 257126 21498 287610 21734
rect 287846 21498 318330 21734
rect 318566 21498 349050 21734
rect 349286 21498 379770 21734
rect 380006 21498 410490 21734
rect 410726 21498 441210 21734
rect 441446 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 471930 21734
rect 472166 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 502650 21734
rect 502886 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 36730 18334
rect 36966 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 67450 18334
rect 67686 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 98170 18334
rect 98406 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 128890 18334
rect 129126 18098 159610 18334
rect 159846 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 190330 18334
rect 190566 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 221050 18334
rect 221286 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 251770 18334
rect 252006 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 282490 18334
rect 282726 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 313210 18334
rect 313446 18098 343930 18334
rect 344166 18098 374650 18334
rect 374886 18098 405370 18334
rect 405606 18098 436090 18334
rect 436326 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 466810 18334
rect 467046 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 497530 18334
rect 497766 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 36730 18014
rect 36966 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 67450 18014
rect 67686 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 98170 18014
rect 98406 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 128890 18014
rect 129126 17778 159610 18014
rect 159846 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 190330 18014
rect 190566 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 221050 18014
rect 221286 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 251770 18014
rect 252006 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 282490 18014
rect 282726 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 313210 18014
rect 313446 17778 343930 18014
rect 344166 17778 374650 18014
rect 374886 17778 405370 18014
rect 405606 17778 436090 18014
rect 436326 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 466810 18014
rect 467046 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 497530 18014
rect 497766 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 31610 14614
rect 31846 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 62330 14614
rect 62566 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 93050 14614
rect 93286 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 123770 14614
rect 124006 14378 154490 14614
rect 154726 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 185210 14614
rect 185446 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 215930 14614
rect 216166 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 246650 14614
rect 246886 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 277370 14614
rect 277606 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 308090 14614
rect 308326 14378 338810 14614
rect 339046 14378 369530 14614
rect 369766 14378 400250 14614
rect 400486 14378 430970 14614
rect 431206 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 461690 14614
rect 461926 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 492410 14614
rect 492646 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 31610 14294
rect 31846 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 62330 14294
rect 62566 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 93050 14294
rect 93286 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 123770 14294
rect 124006 14058 154490 14294
rect 154726 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 185210 14294
rect 185446 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 215930 14294
rect 216166 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 246650 14294
rect 246886 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 277370 14294
rect 277606 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 308090 14294
rect 308326 14058 338810 14294
rect 339046 14058 369530 14294
rect 369766 14058 400250 14294
rect 400486 14058 430970 14294
rect 431206 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 461690 14294
rect 461926 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 492410 14294
rect 492646 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 26490 10894
rect 26726 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 57210 10894
rect 57446 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 87930 10894
rect 88166 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 118650 10894
rect 118886 10658 149370 10894
rect 149606 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 180090 10894
rect 180326 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 210810 10894
rect 211046 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 241530 10894
rect 241766 10658 272250 10894
rect 272486 10658 302970 10894
rect 303206 10658 333690 10894
rect 333926 10658 364410 10894
rect 364646 10658 395130 10894
rect 395366 10658 425850 10894
rect 426086 10658 456570 10894
rect 456806 10658 487290 10894
rect 487526 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 26490 10574
rect 26726 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 57210 10574
rect 57446 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 87930 10574
rect 88166 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 118650 10574
rect 118886 10338 149370 10574
rect 149606 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 180090 10574
rect 180326 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 210810 10574
rect 211046 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 241530 10574
rect 241766 10338 272250 10574
rect 272486 10338 302970 10574
rect 303206 10338 333690 10574
rect 333926 10338 364410 10574
rect 364646 10338 395130 10574
rect 395366 10338 425850 10574
rect 426086 10338 456570 10574
rect 456806 10338 487290 10574
rect 487526 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 21370 7174
rect 21606 6938 52090 7174
rect 52326 6938 82810 7174
rect 83046 6938 113530 7174
rect 113766 6938 144250 7174
rect 144486 6938 174970 7174
rect 175206 6938 205690 7174
rect 205926 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 236410 7174
rect 236646 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 267130 7174
rect 267366 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 297850 7174
rect 298086 6938 328570 7174
rect 328806 6938 359290 7174
rect 359526 6938 390010 7174
rect 390246 6938 420730 7174
rect 420966 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 451450 7174
rect 451686 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 482170 7174
rect 482406 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 21370 6854
rect 21606 6618 52090 6854
rect 52326 6618 82810 6854
rect 83046 6618 113530 6854
rect 113766 6618 144250 6854
rect 144486 6618 174970 6854
rect 175206 6618 205690 6854
rect 205926 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 236410 6854
rect 236646 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 267130 6854
rect 267366 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 297850 6854
rect 298086 6618 328570 6854
rect 328806 6618 359290 6854
rect 359526 6618 390010 6854
rect 390246 6618 420730 6854
rect 420966 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 451450 6854
rect 451686 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 482170 6854
rect 482406 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_IMPACT_HEAD  mprj
timestamp 0
transform 1 0 12000 0 1 3000
box 0 0 500000 600000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 3486 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 584873 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 3486 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 584873 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 602500 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 602500 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 602500 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 602500 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 602500 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 602500 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 2988 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 602500 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 3479 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 584873 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 3479 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 584873 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 3479 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 584873 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 3479 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 584873 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 2988 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 602500 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 2988 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 602500 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 2988 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 602500 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 2988 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 602500 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 602500 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 602500 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 602500 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 602500 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 602500 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 602500 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 2988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 602500 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 3479 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 584873 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 3479 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 584873 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 3479 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 584873 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 3479 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 584873 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 3479 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 584873 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 2988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 602500 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 2988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 602500 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 2988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 602500 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 2988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 602500 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 2988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 602500 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 3479 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 584873 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 3479 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 584873 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 3479 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 584873 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 3479 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 584873 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 3479 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 584873 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 3479 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 584873 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
