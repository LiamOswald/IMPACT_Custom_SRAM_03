** sch_path: /home/impact/Documents/truncation_SRAM/schematic/truncation_SRAM.sch
.subckt truncation_SRAM DataOut0 DataOut1 DataOut2 DataOut3 DataOut4 DataOut5 DataOut6 DataOut7
+ DataOut8 DataOut9 DataOut10 DataOut11 DataOut12 DataOut13 DataOut14 DataOut15 DataOut16 DataOut17 DataOut18
+ DataOut19 DataOut20 DataOut21 DataOut22 DataOut23 DataOut24 DataOut25 DataOut26 DataOut27 DataOut28 DataOut29
+ DataOut30 DataOut31 Trunk0 Trunk1 Trunk2 Trunk3 Trunk4 Trunk5 Trunk6 Trunk7 Trunk8 Trunk9 Trunk10 Trunk11
+ Trunk12 Trunk13 Trunk14 Trunk15 Trunk16 Trunk17 Trunk18 Trunk19 Trunk20 Trunk21 Trunk22 Trunk23 Trunk24
+ Trunk25 Trunk26 Trunk27 Trunk28 Trunk29 Trunk30 Trunk31 DataIn30 DataIn29 DataIn28 DataIn27 DataIn26
+ DataIn25 DataIn24 DataIn23 DataIn22 DataIn21 DataIn20 DataIn19 DataIn18 DataIn17 DataIn16 DataIn15 DataIn14
+ DataIn13 DataIn12 DataIn11 DataIn10 DataIn9 DataIn8 DataIn7 DataIn6 DataIn5 DataIn4 DataIn3 DataIn2 DataIn1
+ DataIn0 DataIn31 PRE writeen readen WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15
+ WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36
+ WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57
+ WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78
+ WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99
+ WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116
+ WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 WL128 WL129 WL130 WL131 WL132 WL133
+ WL134 WL135 WL136 WL137 WL138 WL139 WL140 WL141 WL142 WL143 WL144 WL145 WL146 WL147 WL148 WL149 WL150
+ WL151 WL152 WL153 WL154 WL155 WL156 WL157 WL158 WL159 WL160 WL161 WL162 WL163 WL164 WL165 WL166 WL167
+ WL168 WL169 WL170 WL171 WL172 WL173 WL174 WL175 WL176 WL177 WL178 WL179 WL180 WL181 WL182 WL183 WL184
+ WL185 WL186 WL187 WL188 WL189 WL190 WL191 WL192 WL193 WL194 WL195 WL196 WL197 WL198 WL199 WL200 WL201
+ WL202 WL203 WL204 WL205 WL206 WL207 WL208 WL209 WL210 WL211 WL212 WL213 WL214 WL215 WL216 WL217 WL218
+ WL219 WL220 WL221 WL222 WL223 WL224 WL225 WL226 WL227 WL228 WL229 WL230 WL231 WL232 WL233 WL234 WL235
+ WL236 WL237 WL238 WL239 WL240 WL241 WL242 WL243 WL244 WL245 WL246 WL247 WL248 WL249 WL250 WL251 WL252
+ WL253 WL254 WL255 WL256 WL257 WL258 WL259 WL260 WL261 WL262 WL263 WL264 WL265 WL266 WL267 WL268 WL269
+ WL270 WL271 WL272 WL273 WL274 WL275 WL276 WL277 WL278 WL279 WL280 WL281 WL282 WL283 WL284 WL285 WL286
+ WL287 WL288 WL289 WL290 WL291 WL292 WL293 WL294 WL295 WL296 WL297 WL298 WL299 WL300 WL301 WL302 WL303
+ WL304 WL305 WL306 WL307 WL308 WL309 WL310 WL311 WL312 WL313 WL314 WL315 WL316 WL317 WL318 WL319 WL320
+ WL321 WL322 WL323 WL324 WL325 WL326 WL327 WL328 WL329 WL330 WL331 WL332 WL333 WL334 WL335 WL336 WL337
+ WL338 WL339 WL340 WL341 WL342 WL343 WL344 WL345 WL346 WL347 WL348 WL349 WL350 WL351 WL352 WL353 WL354
+ WL355 WL356 WL357 WL358 WL359 WL360 WL361 WL362 WL363 WL364 WL365 WL366 WL367 WL368 WL369 WL370 WL371
+ WL372 WL373 WL374 WL375 WL376 WL377 WL378 WL379 WL380 WL381 WL382 WL383 WL384 WL385 WL386 WL387 WL388
+ WL389 WL390 WL391 WL392 WL393 WL394 WL395 WL396 WL397 WL398 WL399 WL400 WL401 WL402 WL403 WL404 WL405
+ WL406 WL407 WL408 WL409 WL410 WL411 WL412 WL413 WL414 WL415 WL416 WL417 WL418 WL419 WL420 WL421 WL422
+ WL423 WL424 WL425 WL426 WL427 WL428 WL429 WL430 WL431 WL432 WL433 WL434 WL435 WL436 WL437 WL438 WL439
+ WL440 WL441 WL442 WL443 WL444 WL445 WL446 WL447 WL448 WL449 WL450 WL451 WL452 WL453 WL454 WL455 WL456
+ WL457 WL458 WL459 WL460 WL461 WL462 WL463 WL464 WL465 WL466 WL467 WL468 WL469 WL470 WL471 WL472 WL473
+ WL474 WL475 WL476 WL477 WL478 WL479 WL480 WL481 WL482 WL483 WL484 WL485 WL486 WL487 WL488 WL489 WL490
+ WL491 WL492 WL493 WL494 WL495 WL496 WL497 WL498 WL499 WL500 WL501 WL502 WL503 WL504 WL505 WL506 WL507
+ WL508 WL509 WL510 WL511 WL512 WL513 WL514 WL515 WL516 WL517 WL518 WL519 WL520 WL521 WL522 WL523 WL524
+ WL525 WL526 WL527 WL528 WL529 WL530 WL531 WL532 WL533 WL534 WL535 WL536 WL537 WL538 WL539 WL540 WL541
+ WL542 WL543 WL544 WL545 WL546 WL547 WL548 WL549 WL550 WL551 WL552 WL553 WL554 WL555 WL556 WL557 WL558
+ WL559 WL560 WL561 WL562 WL563 WL564 WL565 WL566 WL567 WL568 WL569 WL570 WL571 WL572 WL573 WL574 WL575
+ WL576 WL577 WL578 WL579 WL580 WL581 WL582 WL583 WL584 WL585 WL586 WL587 WL588 WL589 WL590 WL591 WL592
+ WL593 WL594 WL595 WL596 WL597 WL598 WL599 WL600 WL601 WL602 WL603 WL604 WL605 WL606 WL607 WL608 WL609
+ WL610 WL611 WL612 WL613 WL614 WL615 WL616 WL617 WL618 WL619 WL620 WL621 WL622 WL623 WL624 WL625 WL626
+ WL627 WL628 WL629 WL630 WL631 WL632 WL633 WL634 WL635 WL636 WL637 WL638 WL639 WL640 WL641 WL642 WL643
+ WL644 WL645 WL646 WL647 WL648 WL649 WL650 WL651 WL652 WL653 WL654 WL655 WL656 WL657 WL658 WL659 WL660
+ WL661 WL662 WL663 WL664 WL665 WL666 WL667 WL668 WL669 WL670 WL671 WL672 WL673 WL674 WL675 WL676 WL677
+ WL678 WL679 WL680 WL681 WL682 WL683 WL684 WL685 WL686 WL687 WL688 WL689 WL690 WL691 WL692 WL693 WL694
+ WL695 WL696 WL697 WL698 WL699 WL700 WL701 WL702 WL703 WL704 WL705 WL706 WL707 WL708 WL709 WL710 WL711
+ WL712 WL713 WL714 WL715 WL716 WL717 WL718 WL719 WL720 WL721 WL722 WL723 WL724 WL725 WL726 WL727 WL728
+ WL729 WL730 WL731 WL732 WL733 WL734 WL735 WL736 WL737 WL738 WL739 WL740 WL741 WL742 WL743 WL744 WL745
+ WL746 WL747 WL748 WL749 WL750 WL751 WL752 WL753 WL754 WL755 WL756 WL757 WL758 WL759 WL760 WL761 WL762
+ WL763 WL764 WL765 WL766 WL767 WL768 WL769 WL770 WL771 WL772 WL773 WL774 WL775 WL776 WL777 WL778 WL779
+ WL780 WL781 WL782 WL783 WL784 WL785 WL786 WL787 WL788 WL789 WL790 WL791 WL792 WL793 WL794 WL795 WL796
+ WL797 WL798 WL799 WL800 WL801 WL802 WL803 WL804 WL805 WL806 WL807 WL808 WL809 WL810 WL811 WL812 WL813
+ WL814 WL815 WL816 WL817 WL818 WL819 WL820 WL821 WL822 WL823 WL824 WL825 WL826 WL827 WL828 WL829 WL830
+ WL831 WL832 WL833 WL834 WL835 WL836 WL837 WL838 WL839 WL840 WL841 WL842 WL843 WL844 WL845 WL846 WL847
+ WL848 WL849 WL850 WL851 WL852 WL853 WL854 WL855 WL856 WL857 WL858 WL859 WL860 WL861 WL862 WL863 WL864
+ WL865 WL866 WL867 WL868 WL869 WL870 WL871 WL872 WL873 WL874 WL875 WL876 WL877 WL878 WL879 WL880 WL881
+ WL882 WL883 WL884 WL885 WL886 WL887 WL888 WL889 WL890 WL891 WL892 WL893 WL894 WL895 WL896 WL897 WL898
+ WL899 WL900 WL901 WL902 WL903 WL904 WL905 WL906 WL907 WL908 WL909 WL910 WL911 WL912 WL913 WL914 WL915
+ WL916 WL917 WL918 WL919 WL920 WL921 WL922 WL923 WL924 WL925 WL926 WL927 WL928 WL929 WL930 WL931 WL932
+ WL933 WL934 WL935 WL936 WL937 WL938 WL939 WL940 WL941 WL942 WL943 WL944 WL945 WL946 WL947 WL948 WL949
+ WL950 WL951 WL952 WL953 WL954 WL955 WL956 WL957 WL958 WL959 WL960 WL961 WL962 WL963 WL964 WL965 WL966
+ WL967 WL968 WL969 WL970 WL971 WL972 WL973 WL974 WL975 WL976 WL977 WL978 WL979 WL980 WL981 WL982 WL983
+ WL984 WL985 WL986 WL987 WL988 WL989 WL990 WL991 WL992 WL993 WL994 WL995 WL996 WL997 WL998 WL999 WL1000
+ WL1001 WL1002 WL1003 WL1004 WL1005 WL1006 WL1007 WL1008 WL1009 WL1010 WL1011 WL1012 WL1013 WL1014 WL1015
+ WL1016 WL1017 WL1018 WL1019 WL1020 WL1021 WL1022 WL1023 vssd1 vccd1 Tail_In Byte_Mode_EnableBar
*.PININFO DataOut0:O DataOut1:O DataOut2:O DataOut3:O DataOut4:O DataOut5:O DataOut6:O DataOut7:O
*+ DataOut8:O DataOut9:O DataOut10:O DataOut11:O DataOut12:O DataOut13:O DataOut14:O DataOut15:O DataOut16:O
*+ DataOut17:O DataOut18:O DataOut19:O DataOut20:O DataOut21:O DataOut22:O DataOut23:O DataOut24:O DataOut25:O
*+ DataOut26:O DataOut27:O DataOut28:O DataOut29:O DataOut30:O DataOut31:O Trunk0:I Trunk1:I Trunk2:I Trunk3:I
*+ Trunk4:I Trunk5:I Trunk6:I Trunk7:I Trunk8:I Trunk9:I Trunk10:I Trunk11:I Trunk12:I Trunk13:I Trunk14:I
*+ Trunk15:I Trunk16:I Trunk17:I Trunk18:I Trunk19:I Trunk20:I Trunk21:I Trunk22:I Trunk23:I Trunk24:I Trunk25:I
*+ Trunk26:I Trunk27:I Trunk28:I Trunk29:I Trunk30:I Trunk31:I DataIn30:I DataIn29:I DataIn28:I DataIn27:I
*+ DataIn26:I DataIn25:I DataIn24:I DataIn23:I DataIn22:I DataIn21:I DataIn20:I DataIn19:I DataIn18:I DataIn17:I
*+ DataIn16:I DataIn15:I DataIn14:I DataIn13:I DataIn12:I DataIn11:I DataIn10:I DataIn9:I DataIn8:I DataIn7:I
*+ DataIn6:I DataIn5:I DataIn4:I DataIn3:I DataIn2:I DataIn1:I DataIn0:I DataIn31:I PRE:I writeen:I readen:I
*+ WL0:I WL1:I WL2:I WL3:I WL4:I WL5:I WL6:I WL7:I WL8:I WL9:I WL10:I WL11:I WL12:I WL13:I WL14:I WL15:I
*+ WL16:I WL17:I WL18:I WL19:I WL20:I WL21:I WL22:I WL23:I WL24:I WL25:I WL26:I WL27:I WL28:I WL29:I WL30:I
*+ WL31:I WL32:I WL33:I WL34:I WL35:I WL36:I WL37:I WL38:I WL39:I WL40:I WL41:I WL42:I WL43:I WL44:I WL45:I
*+ WL46:I WL47:I WL48:I WL49:I WL50:I WL51:I WL52:I WL53:I WL54:I WL55:I WL56:I WL57:I WL58:I WL59:I WL60:I
*+ WL61:I WL62:I WL63:I WL64:I WL65:I WL66:I WL67:I WL68:I WL69:I WL70:I WL71:I WL72:I WL73:I WL74:I WL75:I
*+ WL76:I WL77:I WL78:I WL79:I WL80:I WL81:I WL82:I WL83:I WL84:I WL85:I WL86:I WL87:I WL88:I WL89:I WL90:I
*+ WL91:I WL92:I WL93:I WL94:I WL95:I WL96:I WL97:I WL98:I WL99:I WL100:I WL101:I WL102:I WL103:I WL104:I
*+ WL105:I WL106:I WL107:I WL108:I WL109:I WL110:I WL111:I WL112:I WL113:I WL114:I WL115:I WL116:I WL117:I
*+ WL118:I WL119:I WL120:I WL121:I WL122:I WL123:I WL124:I WL125:I WL126:I WL127:I WL128:I WL129:I WL130:I
*+ WL131:I WL132:I WL133:I WL134:I WL135:I WL136:I WL137:I WL138:I WL139:I WL140:I WL141:I WL142:I WL143:I
*+ WL144:I WL145:I WL146:I WL147:I WL148:I WL149:I WL150:I WL151:I WL152:I WL153:I WL154:I WL155:I WL156:I
*+ WL157:I WL158:I WL159:I WL160:I WL161:I WL162:I WL163:I WL164:I WL165:I WL166:I WL167:I WL168:I WL169:I
*+ WL170:I WL171:I WL172:I WL173:I WL174:I WL175:I WL176:I WL177:I WL178:I WL179:I WL180:I WL181:I WL182:I
*+ WL183:I WL184:I WL185:I WL186:I WL187:I WL188:I WL189:I WL190:I WL191:I WL192:I WL193:I WL194:I WL195:I
*+ WL196:I WL197:I WL198:I WL199:I WL200:I WL201:I WL202:I WL203:I WL204:I WL205:I WL206:I WL207:I WL208:I
*+ WL209:I WL210:I WL211:I WL212:I WL213:I WL214:I WL215:I WL216:I WL217:I WL218:I WL219:I WL220:I WL221:I
*+ WL222:I WL223:I WL224:I WL225:I WL226:I WL227:I WL228:I WL229:I WL230:I WL231:I WL232:I WL233:I WL234:I
*+ WL235:I WL236:I WL237:I WL238:I WL239:I WL240:I WL241:I WL242:I WL243:I WL244:I WL245:I WL246:I WL247:I
*+ WL248:I WL249:I WL250:I WL251:I WL252:I WL253:I WL254:I WL255:I WL256:I WL257:I WL258:I WL259:I WL260:I
*+ WL261:I WL262:I WL263:I WL264:I WL265:I WL266:I WL267:I WL268:I WL269:I WL270:I WL271:I WL272:I WL273:I
*+ WL274:I WL275:I WL276:I WL277:I WL278:I WL279:I WL280:I WL281:I WL282:I WL283:I WL284:I WL285:I WL286:I
*+ WL287:I WL288:I WL289:I WL290:I WL291:I WL292:I WL293:I WL294:I WL295:I WL296:I WL297:I WL298:I WL299:I
*+ WL300:I WL301:I WL302:I WL303:I WL304:I WL305:I WL306:I WL307:I WL308:I WL309:I WL310:I WL311:I WL312:I
*+ WL313:I WL314:I WL315:I WL316:I WL317:I WL318:I WL319:I WL320:I WL321:I WL322:I WL323:I WL324:I WL325:I
*+ WL326:I WL327:I WL328:I WL329:I WL330:I WL331:I WL332:I WL333:I WL334:I WL335:I WL336:I WL337:I WL338:I
*+ WL339:I WL340:I WL341:I WL342:I WL343:I WL344:I WL345:I WL346:I WL347:I WL348:I WL349:I WL350:I WL351:I
*+ WL352:I WL353:I WL354:I WL355:I WL356:I WL357:I WL358:I WL359:I WL360:I WL361:I WL362:I WL363:I WL364:I
*+ WL365:I WL366:I WL367:I WL368:I WL369:I WL370:I WL371:I WL372:I WL373:I WL374:I WL375:I WL376:I WL377:I
*+ WL378:I WL379:I WL380:I WL381:I WL382:I WL383:I WL384:I WL385:I WL386:I WL387:I WL388:I WL389:I WL390:I
*+ WL391:I WL392:I WL393:I WL394:I WL395:I WL396:I WL397:I WL398:I WL399:I WL400:I WL401:I WL402:I WL403:I
*+ WL404:I WL405:I WL406:I WL407:I WL408:I WL409:I WL410:I WL411:I WL412:I WL413:I WL414:I WL415:I WL416:I
*+ WL417:I WL418:I WL419:I WL420:I WL421:I WL422:I WL423:I WL424:I WL425:I WL426:I WL427:I WL428:I WL429:I
*+ WL430:I WL431:I WL432:I WL433:I WL434:I WL435:I WL436:I WL437:I WL438:I WL439:I WL440:I WL441:I WL442:I
*+ WL443:I WL444:I WL445:I WL446:I WL447:I WL448:I WL449:I WL450:I WL451:I WL452:I WL453:I WL454:I WL455:I
*+ WL456:I WL457:I WL458:I WL459:I WL460:I WL461:I WL462:I WL463:I WL464:I WL465:I WL466:I WL467:I WL468:I
*+ WL469:I WL470:I WL471:I WL472:I WL473:I WL474:I WL475:I WL476:I WL477:I WL478:I WL479:I WL480:I WL481:I
*+ WL482:I WL483:I WL484:I WL485:I WL486:I WL487:I WL488:I WL489:I WL490:I WL491:I WL492:I WL493:I WL494:I
*+ WL495:I WL496:I WL497:I WL498:I WL499:I WL500:I WL501:I WL502:I WL503:I WL504:I WL505:I WL506:I WL507:I
*+ WL508:I WL509:I WL510:I WL511:I WL512:I WL513:I WL514:I WL515:I WL516:I WL517:I WL518:I WL519:I WL520:I
*+ WL521:I WL522:I WL523:I WL524:I WL525:I WL526:I WL527:I WL528:I WL529:I WL530:I WL531:I WL532:I WL533:I
*+ WL534:I WL535:I WL536:I WL537:I WL538:I WL539:I WL540:I WL541:I WL542:I WL543:I WL544:I WL545:I WL546:I
*+ WL547:I WL548:I WL549:I WL550:I WL551:I WL552:I WL553:I WL554:I WL555:I WL556:I WL557:I WL558:I WL559:I
*+ WL560:I WL561:I WL562:I WL563:I WL564:I WL565:I WL566:I WL567:I WL568:I WL569:I WL570:I WL571:I WL572:I
*+ WL573:I WL574:I WL575:I WL576:I WL577:I WL578:I WL579:I WL580:I WL581:I WL582:I WL583:I WL584:I WL585:I
*+ WL586:I WL587:I WL588:I WL589:I WL590:I WL591:I WL592:I WL593:I WL594:I WL595:I WL596:I WL597:I WL598:I
*+ WL599:I WL600:I WL601:I WL602:I WL603:I WL604:I WL605:I WL606:I WL607:I WL608:I WL609:I WL610:I WL611:I
*+ WL612:I WL613:I WL614:I WL615:I WL616:I WL617:I WL618:I WL619:I WL620:I WL621:I WL622:I WL623:I WL624:I
*+ WL625:I WL626:I WL627:I WL628:I WL629:I WL630:I WL631:I WL632:I WL633:I WL634:I WL635:I WL636:I WL637:I
*+ WL638:I WL639:I WL640:I WL641:I WL642:I WL643:I WL644:I WL645:I WL646:I WL647:I WL648:I WL649:I WL650:I
*+ WL651:I WL652:I WL653:I WL654:I WL655:I WL656:I WL657:I WL658:I WL659:I WL660:I WL661:I WL662:I WL663:I
*+ WL664:I WL665:I WL666:I WL667:I WL668:I WL669:I WL670:I WL671:I WL672:I WL673:I WL674:I WL675:I WL676:I
*+ WL677:I WL678:I WL679:I WL680:I WL681:I WL682:I WL683:I WL684:I WL685:I WL686:I WL687:I WL688:I WL689:I
*+ WL690:I WL691:I WL692:I WL693:I WL694:I WL695:I WL696:I WL697:I WL698:I WL699:I WL700:I WL701:I WL702:I
*+ WL703:I WL704:I WL705:I WL706:I WL707:I WL708:I WL709:I WL710:I WL711:I WL712:I WL713:I WL714:I WL715:I
*+ WL716:I WL717:I WL718:I WL719:I WL720:I WL721:I WL722:I WL723:I WL724:I WL725:I WL726:I WL727:I WL728:I
*+ WL729:I WL730:I WL731:I WL732:I WL733:I WL734:I WL735:I WL736:I WL737:I WL738:I WL739:I WL740:I WL741:I
*+ WL742:I WL743:I WL744:I WL745:I WL746:I WL747:I WL748:I WL749:I WL750:I WL751:I WL752:I WL753:I WL754:I
*+ WL755:I WL756:I WL757:I WL758:I WL759:I WL760:I WL761:I WL762:I WL763:I WL764:I WL765:I WL766:I WL767:I
*+ WL768:I WL769:I WL770:I WL771:I WL772:I WL773:I WL774:I WL775:I WL776:I WL777:I WL778:I WL779:I WL780:I
*+ WL781:I WL782:I WL783:I WL784:I WL785:I WL786:I WL787:I WL788:I WL789:I WL790:I WL791:I WL792:I WL793:I
*+ WL794:I WL795:I WL796:I WL797:I WL798:I WL799:I WL800:I WL801:I WL802:I WL803:I WL804:I WL805:I WL806:I
*+ WL807:I WL808:I WL809:I WL810:I WL811:I WL812:I WL813:I WL814:I WL815:I WL816:I WL817:I WL818:I WL819:I
*+ WL820:I WL821:I WL822:I WL823:I WL824:I WL825:I WL826:I WL827:I WL828:I WL829:I WL830:I WL831:I WL832:I
*+ WL833:I WL834:I WL835:I WL836:I WL837:I WL838:I WL839:I WL840:I WL841:I WL842:I WL843:I WL844:I WL845:I
*+ WL846:I WL847:I WL848:I WL849:I WL850:I WL851:I WL852:I WL853:I WL854:I WL855:I WL856:I WL857:I WL858:I
*+ WL859:I WL860:I WL861:I WL862:I WL863:I WL864:I WL865:I WL866:I WL867:I WL868:I WL869:I WL870:I WL871:I
*+ WL872:I WL873:I WL874:I WL875:I WL876:I WL877:I WL878:I WL879:I WL880:I WL881:I WL882:I WL883:I WL884:I
*+ WL885:I WL886:I WL887:I WL888:I WL889:I WL890:I WL891:I WL892:I WL893:I WL894:I WL895:I WL896:I WL897:I
*+ WL898:I WL899:I WL900:I WL901:I WL902:I WL903:I WL904:I WL905:I WL906:I WL907:I WL908:I WL909:I WL910:I
*+ WL911:I WL912:I WL913:I WL914:I WL915:I WL916:I WL917:I WL918:I WL919:I WL920:I WL921:I WL922:I WL923:I
*+ WL924:I WL925:I WL926:I WL927:I WL928:I WL929:I WL930:I WL931:I WL932:I WL933:I WL934:I WL935:I WL936:I
*+ WL937:I WL938:I WL939:I WL940:I WL941:I WL942:I WL943:I WL944:I WL945:I WL946:I WL947:I WL948:I WL949:I
*+ WL950:I WL951:I WL952:I WL953:I WL954:I WL955:I WL956:I WL957:I WL958:I WL959:I WL960:I WL961:I WL962:I
*+ WL963:I WL964:I WL965:I WL966:I WL967:I WL968:I WL969:I WL970:I WL971:I WL972:I WL973:I WL974:I WL975:I
*+ WL976:I WL977:I WL978:I WL979:I WL980:I WL981:I WL982:I WL983:I WL984:I WL985:I WL986:I WL987:I WL988:I
*+ WL989:I WL990:I WL991:I WL992:I WL993:I WL994:I WL995:I WL996:I WL997:I WL998:I WL999:I WL1000:I WL1001:I
*+ WL1002:I WL1003:I WL1004:I WL1005:I WL1006:I WL1007:I WL1008:I WL1009:I WL1010:I WL1011:I WL1012:I WL1013:I
*+ WL1014:I WL1015:I WL1016:I WL1017:I WL1018:I WL1019:I WL1020:I WL1021:I WL1022:I WL1023:I vssd1:B vccd1:B
*+ Tail_In:I Byte_Mode_EnableBar:B
x1 DataOut31 DataOut30 DataOut29 DataOut28 DataOut27 DataOut26 DataOut25 DataOut24 DataOut23
+ DataOut22 DataOut21 DataOut20 DataOut19 DataOut18 DataOut17 DataOut16 DataOut15 DataOut14 DataOut13 DataOut12
+ DataOut11 DataOut10 DataOut9 DataOut8 DataOut7 DataOut6 DataOut5 DataOut4 DataOut3 DataOut2 DataOut1 DataOut0
+ Trunk0 Trunk1 Trunk2 Trunk3 Trunk4 Trunk5 Trunk6 Trunk7 Trunk8 Trunk9 Trunk10 Trunk11 Trunk12 Trunk13
+ Trunk14 Trunk15 Trunk16 Trunk17 Trunk18 Trunk19 Trunk20 Trunk21 Trunk22 Trunk23 Trunk24 Trunk25 Trunk26
+ Trunk27 Trunk28 Trunk29 Trunk30 Trunk31 Tail_In net1 vccd1 vssd1 Byte_Mode_EnableBar PRE writeen readen
+ DataIn31 DataIn30 DataIn29 DataIn28 DataIn27 DataIn26 DataIn25 DataIn24 DataIn23 DataIn22 DataIn21 DataIn20
+ DataIn19 DataIn18 DataIn17 DataIn16 DataIn15 DataIn14 DataIn13 DataIn12 DataIn11 DataIn10 DataIn9 DataIn8
+ DataIn7 DataIn6 DataIn5 DataIn4 DataIn3 DataIn2 DataIn1 DataIn0 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9
+ WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30
+ WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51
+ WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72
+ WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93
+ WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111
+ WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 WL128
+ WL129 WL130 WL131 WL132 WL133 WL134 WL135 WL136 WL137 WL138 WL139 WL140 WL141 WL142 WL143 WL144 WL145
+ WL146 WL147 WL148 WL149 WL150 WL151 WL152 WL153 WL154 WL155 WL156 WL157 WL158 WL159 WL160 WL161 WL162
+ WL163 WL164 WL165 WL166 WL167 WL168 WL169 WL170 WL171 WL172 WL173 WL174 WL175 WL176 WL177 WL178 WL179
+ WL180 WL181 WL182 WL183 WL184 WL185 WL186 WL187 WL188 WL189 WL190 WL191 WL192 WL193 WL194 WL195 WL196
+ WL197 WL198 WL199 WL200 WL201 WL202 WL203 WL204 WL205 WL206 WL207 WL208 WL209 WL210 WL211 WL212 WL213
+ WL214 WL215 WL216 WL217 WL218 WL219 WL220 WL221 WL222 WL223 WL224 WL225 WL226 WL227 WL228 WL229 WL230
+ WL231 WL232 WL233 WL234 WL235 WL236 WL237 WL238 WL239 WL240 WL241 WL242 WL243 WL244 WL245 WL246 WL247
+ WL248 WL249 WL250 WL251 WL252 WL253 WL254 WL255 WL256 WL257 WL258 WL259 WL260 WL261 WL262 WL263 WL264
+ WL265 WL266 WL267 WL268 WL269 WL270 WL271 WL272 WL273 WL274 WL275 WL276 WL277 WL278 WL279 WL280 WL281
+ WL282 WL283 WL284 WL285 WL286 WL287 WL288 WL289 WL290 WL291 WL292 WL293 WL294 WL295 WL296 WL297 WL298
+ WL299 WL300 WL301 WL302 WL303 WL304 WL305 WL306 WL307 WL308 WL309 WL310 WL311 WL312 WL313 WL314 WL315
+ WL316 WL317 WL318 WL319 WL320 WL321 WL322 WL323 WL324 WL325 WL326 WL327 WL328 WL329 WL330 WL331 WL332
+ WL333 WL334 WL335 WL336 WL337 WL338 WL339 WL340 WL341 WL342 WL343 WL344 WL345 WL346 WL347 WL348 WL349
+ WL350 WL351 WL352 WL353 WL354 WL355 WL356 WL357 WL358 WL359 WL360 WL361 WL362 WL363 WL364 WL365 WL366
+ WL367 WL368 WL369 WL370 WL371 WL372 WL373 WL374 WL375 WL376 WL377 WL378 WL379 WL380 WL381 WL382 WL383
+ WL384 WL385 WL386 WL387 WL388 WL389 WL390 WL391 WL392 WL393 WL394 WL395 WL396 WL397 WL398 WL399 WL400
+ WL401 WL402 WL403 WL404 WL405 WL406 WL407 WL408 WL409 WL410 WL411 WL412 WL413 WL414 WL415 WL416 WL417
+ WL418 WL419 WL420 WL421 WL422 WL423 WL424 WL425 WL426 WL427 WL428 WL429 WL430 WL431 WL432 WL433 WL434
+ WL435 WL436 WL437 WL438 WL439 WL440 WL441 WL442 WL443 WL444 WL445 WL446 WL447 WL448 WL449 WL450 WL451
+ WL452 WL453 WL454 WL455 WL456 WL457 WL458 WL459 WL460 WL461 WL462 WL463 WL464 WL465 WL466 WL467 WL468
+ WL469 WL470 WL471 WL472 WL473 WL474 WL475 WL476 WL477 WL478 WL479 WL480 WL481 WL482 WL483 WL484 WL485
+ WL486 WL487 WL488 WL489 WL490 WL491 WL492 WL493 WL494 WL495 WL496 WL497 WL498 WL499 WL500 WL501 WL502
+ WL503 WL504 WL505 WL506 WL507 WL508 WL509 WL510 WL511 WL512 WL513 WL514 WL515 WL516 WL517 WL518 WL519
+ WL520 WL521 WL522 WL523 WL524 WL525 WL526 WL527 WL528 WL529 WL530 WL531 WL532 WL533 WL534 WL535 WL536
+ WL537 WL538 WL539 WL540 WL541 WL542 WL543 WL544 WL545 WL546 WL547 WL548 WL549 WL550 WL551 WL552 WL553
+ WL554 WL555 WL556 WL557 WL558 WL559 WL560 WL561 WL562 WL563 WL564 WL565 WL566 WL567 WL568 WL569 WL570
+ WL571 WL572 WL573 WL574 WL575 WL576 WL577 WL578 WL579 WL580 WL581 WL582 WL583 WL584 WL585 WL586 WL587
+ WL588 WL589 WL590 WL591 WL592 WL593 WL594 WL595 WL596 WL597 WL598 WL599 WL600 WL601 WL602 WL603 WL604
+ WL605 WL606 WL607 WL608 WL609 WL610 WL611 WL612 WL613 WL614 WL615 WL616 WL617 WL618 WL619 WL620 WL621
+ WL622 WL623 WL624 WL625 WL626 WL627 WL628 WL629 WL630 WL631 WL632 WL633 WL634 WL635 WL636 WL637 WL638
+ WL639 WL640 WL641 WL642 WL643 WL644 WL645 WL646 WL647 WL648 WL649 WL650 WL651 WL652 WL653 WL654 WL655
+ WL656 WL657 WL658 WL659 WL660 WL661 WL662 WL663 WL664 WL665 WL666 WL667 WL668 WL669 WL670 WL671 WL672
+ WL673 WL674 WL675 WL676 WL677 WL678 WL679 WL680 WL681 WL682 WL683 WL684 WL685 WL686 WL687 WL688 WL689
+ WL690 WL691 WL692 WL693 WL694 WL695 WL696 WL697 WL698 WL699 WL700 WL701 WL702 WL703 WL704 WL705 WL706
+ WL707 WL708 WL709 WL710 WL711 WL712 WL713 WL714 WL715 WL716 WL717 WL718 WL719 WL720 WL721 WL722 WL723
+ WL724 WL725 WL726 WL727 WL728 WL729 WL730 WL731 WL732 WL733 WL734 WL735 WL736 WL737 WL738 WL739 WL740
+ WL741 WL742 WL743 WL744 WL745 WL746 WL747 WL748 WL749 WL750 WL751 WL752 WL753 WL754 WL755 WL756 WL757
+ WL758 WL759 WL760 WL761 WL762 WL763 WL764 WL765 WL766 WL767 WL768 WL769 WL770 WL771 WL772 WL773 WL774
+ WL775 WL776 WL777 WL778 WL779 WL780 WL781 WL782 WL783 WL784 WL785 WL786 WL787 WL788 WL789 WL790 WL791
+ WL792 WL793 WL794 WL795 WL796 WL797 WL798 WL799 WL800 WL801 WL802 WL803 WL804 WL805 WL806 WL807 WL808
+ WL809 WL810 WL811 WL812 WL813 WL814 WL815 WL816 WL817 WL818 WL819 WL820 WL821 WL822 WL823 WL824 WL825
+ WL826 WL827 WL828 WL829 WL830 WL831 WL832 WL833 WL834 WL835 WL836 WL837 WL838 WL839 WL840 WL841 WL842
+ WL843 WL844 WL845 WL846 WL847 WL848 WL849 WL850 WL851 WL852 WL853 WL854 WL855 WL856 WL857 WL858 WL859
+ WL860 WL861 WL862 WL863 WL864 WL865 WL866 WL867 WL868 WL869 WL870 WL871 WL872 WL873 WL874 WL875 WL876
+ WL877 WL878 WL879 WL880 WL881 WL882 WL883 WL884 WL885 WL886 WL887 WL888 WL889 WL890 WL891 WL892 WL893
+ WL894 WL895 WL896 WL897 WL898 WL899 WL900 WL901 WL902 WL903 WL904 WL905 WL906 WL907 WL908 WL909 WL910
+ WL911 WL912 WL913 WL914 WL915 WL916 WL917 WL918 WL919 WL920 WL921 WL922 WL923 WL924 WL925 WL926 WL927
+ WL928 WL929 WL930 WL931 WL932 WL933 WL934 WL935 WL936 WL937 WL938 WL939 WL940 WL941 WL942 WL943 WL944
+ WL945 WL946 WL947 WL948 WL949 WL950 WL951 WL952 WL953 WL954 WL955 WL956 WL957 WL958 WL959 WL960 WL961
+ WL962 WL963 WL964 WL965 WL966 WL967 WL968 WL969 WL970 WL971 WL972 WL973 WL974 WL975 WL976 WL977 WL978
+ WL979 WL980 WL981 WL982 WL983 WL984 WL985 WL986 WL987 WL988 WL989 WL990 WL991 WL992 WL993 WL994 WL995
+ WL996 WL997 WL998 WL999 WL1000 WL1001 WL1002 WL1003 WL1004 WL1005 WL1006 WL1007 WL1008 WL1009 WL1010
+ WL1011 WL1012 WL1013 WL1014 WL1015 WL1016 WL1017 WL1018 WL1019 WL1020 WL1021 WL1022 WL1023
+ 32x1024_truncation_memory
.ends

* expanding   symbol:
*+  /home/impact/Documents/truncation_SRAM/schematic/32x1024_truncation_memory.sym # of pins=1128
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/32x1024_truncation_memory.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/32x1024_truncation_memory.sch
.subckt 32x1024_truncation_memory DataOut31 DataOut30 DataOut29 DataOut28 DataOut27 DataOut26
+ DataOut25 DataOut24 DataOut23 DataOut22 DataOut21 DataOut20 DataOut19 DataOut18 DataOut17 DataOut16 DataOut15
+ DataOut14 DataOut13 DataOut12 DataOut11 DataOut10 DataOut9 DataOut8 DataOut7 DataOut6 DataOut5 DataOut4
+ DataOut3 DataOut2 DataOut1 DataOut0 Trunk0 Trunk1 Trunk2 Trunk3 Trunk4 Trunk5 Trunk6 Trunk7 Trunk8 Trunk9
+ Trunk10 Trunk11 Trunk12 Trunk13 Trunk14 Trunk15 Trunk16 Trunk17 Trunk18 Trunk19 Trunk20 Trunk21 Trunk22
+ Trunk23 Trunk24 Trunk25 Trunk26 Trunk27 Trunk28 Trunk29 Trunk30 Trunk31 Tail_In Tail_Out vccd1 vssd1
+ Byte_Mode_EnableBar PRE writeen readen DataIn31 DataIn30 DataIn29 DataIn28 DataIn27 DataIn26 DataIn25 DataIn24 DataIn23
+ DataIn22 DataIn21 DataIn20 DataIn19 DataIn18 DataIn17 DataIn16 DataIn15 DataIn14 DataIn13 DataIn12 DataIn11
+ DataIn10 DataIn9 DataIn8 DataIn7 DataIn6 DataIn5 DataIn4 DataIn3 DataIn2 DataIn1 DataIn0 WL0 WL1 WL2 WL3 WL4
+ WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25
+ WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46
+ WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67
+ WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88
+ WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107
+ WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124
+ WL125 WL126 WL127 WL128 WL129 WL130 WL131 WL132 WL133 WL134 WL135 WL136 WL137 WL138 WL139 WL140 WL141
+ WL142 WL143 WL144 WL145 WL146 WL147 WL148 WL149 WL150 WL151 WL152 WL153 WL154 WL155 WL156 WL157 WL158
+ WL159 WL160 WL161 WL162 WL163 WL164 WL165 WL166 WL167 WL168 WL169 WL170 WL171 WL172 WL173 WL174 WL175
+ WL176 WL177 WL178 WL179 WL180 WL181 WL182 WL183 WL184 WL185 WL186 WL187 WL188 WL189 WL190 WL191 WL192
+ WL193 WL194 WL195 WL196 WL197 WL198 WL199 WL200 WL201 WL202 WL203 WL204 WL205 WL206 WL207 WL208 WL209
+ WL210 WL211 WL212 WL213 WL214 WL215 WL216 WL217 WL218 WL219 WL220 WL221 WL222 WL223 WL224 WL225 WL226
+ WL227 WL228 WL229 WL230 WL231 WL232 WL233 WL234 WL235 WL236 WL237 WL238 WL239 WL240 WL241 WL242 WL243
+ WL244 WL245 WL246 WL247 WL248 WL249 WL250 WL251 WL252 WL253 WL254 WL255 WL256 WL257 WL258 WL259 WL260
+ WL261 WL262 WL263 WL264 WL265 WL266 WL267 WL268 WL269 WL270 WL271 WL272 WL273 WL274 WL275 WL276 WL277
+ WL278 WL279 WL280 WL281 WL282 WL283 WL284 WL285 WL286 WL287 WL288 WL289 WL290 WL291 WL292 WL293 WL294
+ WL295 WL296 WL297 WL298 WL299 WL300 WL301 WL302 WL303 WL304 WL305 WL306 WL307 WL308 WL309 WL310 WL311
+ WL312 WL313 WL314 WL315 WL316 WL317 WL318 WL319 WL320 WL321 WL322 WL323 WL324 WL325 WL326 WL327 WL328
+ WL329 WL330 WL331 WL332 WL333 WL334 WL335 WL336 WL337 WL338 WL339 WL340 WL341 WL342 WL343 WL344 WL345
+ WL346 WL347 WL348 WL349 WL350 WL351 WL352 WL353 WL354 WL355 WL356 WL357 WL358 WL359 WL360 WL361 WL362
+ WL363 WL364 WL365 WL366 WL367 WL368 WL369 WL370 WL371 WL372 WL373 WL374 WL375 WL376 WL377 WL378 WL379
+ WL380 WL381 WL382 WL383 WL384 WL385 WL386 WL387 WL388 WL389 WL390 WL391 WL392 WL393 WL394 WL395 WL396
+ WL397 WL398 WL399 WL400 WL401 WL402 WL403 WL404 WL405 WL406 WL407 WL408 WL409 WL410 WL411 WL412 WL413
+ WL414 WL415 WL416 WL417 WL418 WL419 WL420 WL421 WL422 WL423 WL424 WL425 WL426 WL427 WL428 WL429 WL430
+ WL431 WL432 WL433 WL434 WL435 WL436 WL437 WL438 WL439 WL440 WL441 WL442 WL443 WL444 WL445 WL446 WL447
+ WL448 WL449 WL450 WL451 WL452 WL453 WL454 WL455 WL456 WL457 WL458 WL459 WL460 WL461 WL462 WL463 WL464
+ WL465 WL466 WL467 WL468 WL469 WL470 WL471 WL472 WL473 WL474 WL475 WL476 WL477 WL478 WL479 WL480 WL481
+ WL482 WL483 WL484 WL485 WL486 WL487 WL488 WL489 WL490 WL491 WL492 WL493 WL494 WL495 WL496 WL497 WL498
+ WL499 WL500 WL501 WL502 WL503 WL504 WL505 WL506 WL507 WL508 WL509 WL510 WL511 WL512 WL513 WL514 WL515
+ WL516 WL517 WL518 WL519 WL520 WL521 WL522 WL523 WL524 WL525 WL526 WL527 WL528 WL529 WL530 WL531 WL532
+ WL533 WL534 WL535 WL536 WL537 WL538 WL539 WL540 WL541 WL542 WL543 WL544 WL545 WL546 WL547 WL548 WL549
+ WL550 WL551 WL552 WL553 WL554 WL555 WL556 WL557 WL558 WL559 WL560 WL561 WL562 WL563 WL564 WL565 WL566
+ WL567 WL568 WL569 WL570 WL571 WL572 WL573 WL574 WL575 WL576 WL577 WL578 WL579 WL580 WL581 WL582 WL583
+ WL584 WL585 WL586 WL587 WL588 WL589 WL590 WL591 WL592 WL593 WL594 WL595 WL596 WL597 WL598 WL599 WL600
+ WL601 WL602 WL603 WL604 WL605 WL606 WL607 WL608 WL609 WL610 WL611 WL612 WL613 WL614 WL615 WL616 WL617
+ WL618 WL619 WL620 WL621 WL622 WL623 WL624 WL625 WL626 WL627 WL628 WL629 WL630 WL631 WL632 WL633 WL634
+ WL635 WL636 WL637 WL638 WL639 WL640 WL641 WL642 WL643 WL644 WL645 WL646 WL647 WL648 WL649 WL650 WL651
+ WL652 WL653 WL654 WL655 WL656 WL657 WL658 WL659 WL660 WL661 WL662 WL663 WL664 WL665 WL666 WL667 WL668
+ WL669 WL670 WL671 WL672 WL673 WL674 WL675 WL676 WL677 WL678 WL679 WL680 WL681 WL682 WL683 WL684 WL685
+ WL686 WL687 WL688 WL689 WL690 WL691 WL692 WL693 WL694 WL695 WL696 WL697 WL698 WL699 WL700 WL701 WL702
+ WL703 WL704 WL705 WL706 WL707 WL708 WL709 WL710 WL711 WL712 WL713 WL714 WL715 WL716 WL717 WL718 WL719
+ WL720 WL721 WL722 WL723 WL724 WL725 WL726 WL727 WL728 WL729 WL730 WL731 WL732 WL733 WL734 WL735 WL736
+ WL737 WL738 WL739 WL740 WL741 WL742 WL743 WL744 WL745 WL746 WL747 WL748 WL749 WL750 WL751 WL752 WL753
+ WL754 WL755 WL756 WL757 WL758 WL759 WL760 WL761 WL762 WL763 WL764 WL765 WL766 WL767 WL768 WL769 WL770
+ WL771 WL772 WL773 WL774 WL775 WL776 WL777 WL778 WL779 WL780 WL781 WL782 WL783 WL784 WL785 WL786 WL787
+ WL788 WL789 WL790 WL791 WL792 WL793 WL794 WL795 WL796 WL797 WL798 WL799 WL800 WL801 WL802 WL803 WL804
+ WL805 WL806 WL807 WL808 WL809 WL810 WL811 WL812 WL813 WL814 WL815 WL816 WL817 WL818 WL819 WL820 WL821
+ WL822 WL823 WL824 WL825 WL826 WL827 WL828 WL829 WL830 WL831 WL832 WL833 WL834 WL835 WL836 WL837 WL838
+ WL839 WL840 WL841 WL842 WL843 WL844 WL845 WL846 WL847 WL848 WL849 WL850 WL851 WL852 WL853 WL854 WL855
+ WL856 WL857 WL858 WL859 WL860 WL861 WL862 WL863 WL864 WL865 WL866 WL867 WL868 WL869 WL870 WL871 WL872
+ WL873 WL874 WL875 WL876 WL877 WL878 WL879 WL880 WL881 WL882 WL883 WL884 WL885 WL886 WL887 WL888 WL889
+ WL890 WL891 WL892 WL893 WL894 WL895 WL896 WL897 WL898 WL899 WL900 WL901 WL902 WL903 WL904 WL905 WL906
+ WL907 WL908 WL909 WL910 WL911 WL912 WL913 WL914 WL915 WL916 WL917 WL918 WL919 WL920 WL921 WL922 WL923
+ WL924 WL925 WL926 WL927 WL928 WL929 WL930 WL931 WL932 WL933 WL934 WL935 WL936 WL937 WL938 WL939 WL940
+ WL941 WL942 WL943 WL944 WL945 WL946 WL947 WL948 WL949 WL950 WL951 WL952 WL953 WL954 WL955 WL956 WL957
+ WL958 WL959 WL960 WL961 WL962 WL963 WL964 WL965 WL966 WL967 WL968 WL969 WL970 WL971 WL972 WL973 WL974
+ WL975 WL976 WL977 WL978 WL979 WL980 WL981 WL982 WL983 WL984 WL985 WL986 WL987 WL988 WL989 WL990 WL991
+ WL992 WL993 WL994 WL995 WL996 WL997 WL998 WL999 WL1000 WL1001 WL1002 WL1003 WL1004 WL1005 WL1006 WL1007
+ WL1008 WL1009 WL1010 WL1011 WL1012 WL1013 WL1014 WL1015 WL1016 WL1017 WL1018 WL1019 WL1020 WL1021 WL1022
+ WL1023
*.PININFO vssd1:B vccd1:B WL0:I WL1:I WL2:I WL3:I WL4:I WL5:I WL6:I WL7:I WL8:I WL9:I WL10:I WL11:I
*+ WL12:I WL13:I WL14:I WL15:I WL16:I WL17:I WL18:I WL19:I WL20:I WL21:I WL22:I WL23:I WL24:I WL25:I WL26:I
*+ WL27:I WL28:I WL29:I WL30:I WL31:I WL32:I WL33:I WL34:I WL35:I WL36:I WL37:I WL38:I WL39:I WL40:I WL41:I
*+ WL42:I WL43:I WL44:I WL45:I WL46:I WL47:I WL48:I WL49:I WL50:I WL51:I WL52:I WL53:I WL54:I WL55:I WL56:I
*+ WL57:I WL58:I WL59:I WL60:I WL61:I WL62:I WL63:I WL64:I WL65:I WL66:I WL67:I WL68:I WL69:I WL70:I WL71:I
*+ WL72:I WL73:I WL74:I WL75:I WL76:I WL77:I WL78:I WL79:I WL80:I WL81:I WL82:I WL83:I WL84:I WL85:I WL86:I
*+ WL87:I WL88:I WL89:I WL90:I WL91:I WL92:I WL93:I WL94:I WL95:I WL96:I WL97:I WL98:I WL99:I WL100:I WL101:I
*+ WL102:I WL103:I WL104:I WL105:I WL106:I WL107:I WL108:I WL109:I WL110:I WL111:I WL112:I WL113:I WL114:I
*+ WL115:I WL116:I WL117:I WL118:I WL119:I WL120:I WL121:I WL122:I WL123:I WL124:I WL125:I WL126:I WL127:I
*+ WL128:I WL129:I WL130:I WL131:I WL132:I WL133:I WL134:I WL135:I WL136:I WL137:I WL138:I WL139:I WL140:I
*+ WL141:I WL142:I WL143:I WL144:I WL145:I WL146:I WL147:I WL148:I WL149:I WL150:I WL151:I WL152:I WL153:I
*+ WL154:I WL155:I WL156:I WL157:I WL158:I WL159:I WL160:I WL161:I WL162:I WL163:I WL164:I WL165:I WL166:I
*+ WL167:I WL168:I WL169:I WL170:I WL171:I WL172:I WL173:I WL174:I WL175:I WL176:I WL177:I WL178:I WL179:I
*+ WL180:I WL181:I WL182:I WL183:I WL184:I WL185:I WL186:I WL187:I WL188:I WL189:I WL190:I WL191:I WL192:I
*+ WL193:I WL194:I WL195:I WL196:I WL197:I WL198:I WL199:I WL200:I WL201:I WL202:I WL203:I WL204:I WL205:I
*+ WL206:I WL207:I WL208:I WL209:I WL210:I WL211:I WL212:I WL213:I WL214:I WL215:I WL216:I WL217:I WL218:I
*+ WL219:I WL220:I WL221:I WL222:I WL223:I WL224:I WL225:I WL226:I WL227:I WL228:I WL229:I WL230:I WL231:I
*+ WL232:I WL233:I WL234:I WL235:I WL236:I WL237:I WL238:I WL239:I WL240:I WL241:I WL242:I WL243:I WL244:I
*+ WL245:I WL246:I WL247:I WL248:I WL249:I WL250:I WL251:I WL252:I WL253:I WL254:I WL255:I WL256:I WL257:I
*+ WL258:I WL259:I WL260:I WL261:I WL262:I WL263:I WL264:I WL265:I WL266:I WL267:I WL268:I WL269:I WL270:I
*+ WL271:I WL272:I WL273:I WL274:I WL275:I WL276:I WL277:I WL278:I WL279:I WL280:I WL281:I WL282:I WL283:I
*+ WL284:I WL285:I WL286:I WL287:I WL288:I WL289:I WL290:I WL291:I WL292:I WL293:I WL294:I WL295:I WL296:I
*+ WL297:I WL298:I WL299:I WL300:I WL301:I WL302:I WL303:I WL304:I WL305:I WL306:I WL307:I WL308:I WL309:I
*+ WL310:I WL311:I WL312:I WL313:I WL314:I WL315:I WL316:I WL317:I WL318:I WL319:I WL320:I WL321:I WL322:I
*+ WL323:I WL324:I WL325:I WL326:I WL327:I WL328:I WL329:I WL330:I WL331:I WL332:I WL333:I WL334:I WL335:I
*+ WL336:I WL337:I WL338:I WL339:I WL340:I WL341:I WL342:I WL343:I WL344:I WL345:I WL346:I WL347:I WL348:I
*+ WL349:I WL350:I WL351:I WL352:I WL353:I WL354:I WL355:I WL356:I WL357:I WL358:I WL359:I WL360:I WL361:I
*+ WL362:I WL363:I WL364:I WL365:I WL366:I WL367:I WL368:I WL369:I WL370:I WL371:I WL372:I WL373:I WL374:I
*+ WL375:I WL376:I WL377:I WL378:I WL379:I WL380:I WL381:I WL382:I WL383:I WL384:I WL385:I WL386:I WL387:I
*+ WL388:I WL389:I WL390:I WL391:I WL392:I WL393:I WL394:I WL395:I WL396:I WL397:I WL398:I WL399:I WL400:I
*+ WL401:I WL402:I WL403:I WL404:I WL405:I WL406:I WL407:I WL408:I WL409:I WL410:I WL411:I WL412:I WL413:I
*+ WL414:I WL415:I WL416:I WL417:I WL418:I WL419:I WL420:I WL421:I WL422:I WL423:I WL424:I WL425:I WL426:I
*+ WL427:I WL428:I WL429:I WL430:I WL431:I WL432:I WL433:I WL434:I WL435:I WL436:I WL437:I WL438:I WL439:I
*+ WL440:I WL441:I WL442:I WL443:I WL444:I WL445:I WL446:I WL447:I WL448:I WL449:I WL450:I WL451:I WL452:I
*+ WL453:I WL454:I WL455:I WL456:I WL457:I WL458:I WL459:I WL460:I WL461:I WL462:I WL463:I WL464:I WL465:I
*+ WL466:I WL467:I WL468:I WL469:I WL470:I WL471:I WL472:I WL473:I WL474:I WL475:I WL476:I WL477:I WL478:I
*+ WL479:I WL480:I WL481:I WL482:I WL483:I WL484:I WL485:I WL486:I WL487:I WL488:I WL489:I WL490:I WL491:I
*+ WL492:I WL493:I WL494:I WL495:I WL496:I WL497:I WL498:I WL499:I WL500:I WL501:I WL502:I WL503:I WL504:I
*+ WL505:I WL506:I WL507:I WL508:I WL509:I WL510:I WL511:I WL512:I WL513:I WL514:I WL515:I WL516:I WL517:I
*+ WL518:I WL519:I WL520:I WL521:I WL522:I WL523:I WL524:I WL525:I WL526:I WL527:I WL528:I WL529:I WL530:I
*+ WL531:I WL532:I WL533:I WL534:I WL535:I WL536:I WL537:I WL538:I WL539:I WL540:I WL541:I WL542:I WL543:I
*+ WL544:I WL545:I WL546:I WL547:I WL548:I WL549:I WL550:I WL551:I WL552:I WL553:I WL554:I WL555:I WL556:I
*+ WL557:I WL558:I WL559:I WL560:I WL561:I WL562:I WL563:I WL564:I WL565:I WL566:I WL567:I WL568:I WL569:I
*+ WL570:I WL571:I WL572:I WL573:I WL574:I WL575:I WL576:I WL577:I WL578:I WL579:I WL580:I WL581:I WL582:I
*+ WL583:I WL584:I WL585:I WL586:I WL587:I WL588:I WL589:I WL590:I WL591:I WL592:I WL593:I WL594:I WL595:I
*+ WL596:I WL597:I WL598:I WL599:I WL600:I WL601:I WL602:I WL603:I WL604:I WL605:I WL606:I WL607:I WL608:I
*+ WL609:I WL610:I WL611:I WL612:I WL613:I WL614:I WL615:I WL616:I WL617:I WL618:I WL619:I WL620:I WL621:I
*+ WL622:I WL623:I WL624:I WL625:I WL626:I WL627:I WL628:I WL629:I WL630:I WL631:I WL632:I WL633:I WL634:I
*+ WL635:I WL636:I WL637:I WL638:I WL639:I WL640:I WL641:I WL642:I WL643:I WL644:I WL645:I WL646:I WL647:I
*+ WL648:I WL649:I WL650:I WL651:I WL652:I WL653:I WL654:I WL655:I WL656:I WL657:I WL658:I WL659:I WL660:I
*+ WL661:I WL662:I WL663:I WL664:I WL665:I WL666:I WL667:I WL668:I WL669:I WL670:I WL671:I WL672:I WL673:I
*+ WL674:I WL675:I WL676:I WL677:I WL678:I WL679:I WL680:I WL681:I WL682:I WL683:I WL684:I WL685:I WL686:I
*+ WL687:I WL688:I WL689:I WL690:I WL691:I WL692:I WL693:I WL694:I WL695:I WL696:I WL697:I WL698:I WL699:I
*+ WL700:I WL701:I WL702:I WL703:I WL704:I WL705:I WL706:I WL707:I WL708:I WL709:I WL710:I WL711:I WL712:I
*+ WL713:I WL714:I WL715:I WL716:I WL717:I WL718:I WL719:I WL720:I WL721:I WL722:I WL723:I WL724:I WL725:I
*+ WL726:I WL727:I WL728:I WL729:I WL730:I WL731:I WL732:I WL733:I WL734:I WL735:I WL736:I WL737:I WL738:I
*+ WL739:I WL740:I WL741:I WL742:I WL743:I WL744:I WL745:I WL746:I WL747:I WL748:I WL749:I WL750:I WL751:I
*+ WL752:I WL753:I WL754:I WL755:I WL756:I WL757:I WL758:I WL759:I WL760:I WL761:I WL762:I WL763:I WL764:I
*+ WL765:I WL766:I WL767:I WL768:I WL769:I WL770:I WL771:I WL772:I WL773:I WL774:I WL775:I WL776:I WL777:I
*+ WL778:I WL779:I WL780:I WL781:I WL782:I WL783:I WL784:I WL785:I WL786:I WL787:I WL788:I WL789:I WL790:I
*+ WL791:I WL792:I WL793:I WL794:I WL795:I WL796:I WL797:I WL798:I WL799:I WL800:I WL801:I WL802:I WL803:I
*+ WL804:I WL805:I WL806:I WL807:I WL808:I WL809:I WL810:I WL811:I WL812:I WL813:I WL814:I WL815:I WL816:I
*+ WL817:I WL818:I WL819:I WL820:I WL821:I WL822:I WL823:I WL824:I WL825:I WL826:I WL827:I WL828:I WL829:I
*+ WL830:I WL831:I WL832:I WL833:I WL834:I WL835:I WL836:I WL837:I WL838:I WL839:I WL840:I WL841:I WL842:I
*+ WL843:I WL844:I WL845:I WL846:I WL847:I WL848:I WL849:I WL850:I WL851:I WL852:I WL853:I WL854:I WL855:I
*+ WL856:I WL857:I WL858:I WL859:I WL860:I WL861:I WL862:I WL863:I WL864:I WL865:I WL866:I WL867:I WL868:I
*+ WL869:I WL870:I WL871:I WL872:I WL873:I WL874:I WL875:I WL876:I WL877:I WL878:I WL879:I WL880:I WL881:I
*+ WL882:I WL883:I WL884:I WL885:I WL886:I WL887:I WL888:I WL889:I WL890:I WL891:I WL892:I WL893:I WL894:I
*+ WL895:I WL896:I WL897:I WL898:I WL899:I WL900:I WL901:I WL902:I WL903:I WL904:I WL905:I WL906:I WL907:I
*+ WL908:I WL909:I WL910:I WL911:I WL912:I WL913:I WL914:I WL915:I WL916:I WL917:I WL918:I WL919:I WL920:I
*+ WL921:I WL922:I WL923:I WL924:I WL925:I WL926:I WL927:I WL928:I WL929:I WL930:I WL931:I WL932:I WL933:I
*+ WL934:I WL935:I WL936:I WL937:I WL938:I WL939:I WL940:I WL941:I WL942:I WL943:I WL944:I WL945:I WL946:I
*+ WL947:I WL948:I WL949:I WL950:I WL951:I WL952:I WL953:I WL954:I WL955:I WL956:I WL957:I WL958:I WL959:I
*+ WL960:I WL961:I WL962:I WL963:I WL964:I WL965:I WL966:I WL967:I WL968:I WL969:I WL970:I WL971:I WL972:I
*+ WL973:I WL974:I WL975:I WL976:I WL977:I WL978:I WL979:I WL980:I WL981:I WL982:I WL983:I WL984:I WL985:I
*+ WL986:I WL987:I WL988:I WL989:I WL990:I WL991:I WL992:I WL993:I WL994:I WL995:I WL996:I WL997:I WL998:I
*+ WL999:I WL1000:I WL1001:I WL1002:I WL1003:I WL1004:I WL1005:I WL1006:I WL1007:I WL1008:I WL1009:I WL1010:I
*+ WL1011:I WL1012:I WL1013:I WL1014:I WL1015:I WL1016:I WL1017:I WL1018:I WL1019:I WL1020:I WL1021:I WL1022:I
*+ WL1023:I DataIn30:I DataIn29:I DataIn28:I DataIn27:I DataIn26:I DataIn25:I DataIn24:I DataIn23:I DataIn22:I
*+ DataIn21:I DataIn20:I DataIn19:I DataIn18:I DataIn17:I DataIn16:I DataIn15:I DataIn14:I DataIn13:I DataIn12:I
*+ DataIn11:I DataIn10:I DataIn9:I DataIn8:I DataIn7:I DataIn6:I DataIn5:I DataIn4:I DataIn3:I DataIn2:I
*+ DataIn1:I DataIn0:I DataIn31:I PRE:I writeen:I readen:I Trunk0:I Trunk1:I Trunk2:I Trunk3:I Trunk4:I Trunk5:I
*+ Trunk6:I Trunk7:I Trunk8:I Trunk9:I Trunk10:I Trunk11:I Trunk12:I Trunk13:I Trunk14:I Trunk15:I Trunk16:I
*+ Trunk17:I Trunk18:I Trunk19:I Trunk20:I Trunk21:I Trunk22:I Trunk23:I Trunk24:I Trunk25:I Trunk26:I Trunk27:I
*+ Trunk28:I Trunk29:I Trunk30:I Trunk31:I Tail_In:I Byte_Mode_EnableBar:B Tail_Out:O DataOut0:O DataOut1:O
*+ DataOut2:O DataOut3:O DataOut4:O DataOut5:O DataOut6:O DataOut7:O DataOut8:O DataOut9:O DataOut10:O
*+ DataOut11:O DataOut12:O DataOut13:O DataOut14:O DataOut15:O DataOut16:O DataOut17:O DataOut18:O DataOut19:O
*+ DataOut20:O DataOut21:O DataOut22:O DataOut23:O DataOut24:O DataOut25:O DataOut26:O DataOut27:O DataOut28:O
*+ DataOut29:O DataOut30:O DataOut31:O
x1 vccd1 net38 net39 net40 net41 net42 net43 net44 net45 net46 net47 net48 net49 net50 net51 net52
+ net53 net2 net1 net4 net3 net6 net5 net8 net7 net10 net9 net12 net11 net14 net13 net16 net15 net18 net17
+ net20 net19 net22 net21 net24 net23 net26 net25 net28 net27 net30 net29 net32 net31 net54 net34 net33
+ net36 net35 net37 net55 net56 net57 net58 net59 net60 net61 net62 net63 net64 vssd1 PRE writeen readen
+ DataIn31 DataIn30 DataIn29 DataIn28 DataIn27 DataIn26 DataIn25 DataIn24 DataIn23 DataIn22 DataIn21 DataIn20
+ DataIn19 DataIn18 DataIn17 DataIn16 DataIn15 DataIn14 DataIn13 DataIn12 DataIn11 DataIn10 DataIn9 DataIn8
+ DataIn7 DataIn6 DataIn5 DataIn4 DataIn3 DataIn2 DataIn1 DataIn0 Read31 Read30 Read29 Read28 Read27 Read26
+ Read25 Read24 Read23 Read22 Read21 Read20 Read19 Read18 Read17 Read16 Read15 Read14 Read13 Read12 Read11
+ Read10 Read9 Read8 Read7 Read6 Read5 Read4 Read3 Read2 Read1 Read0 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9
+ WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30
+ WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51
+ WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72
+ WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93
+ WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111
+ WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 WL128
+ WL129 WL130 WL131 WL132 WL133 WL134 WL135 WL136 WL137 WL138 WL139 WL140 WL141 WL142 WL143 WL144 WL145
+ WL146 WL147 WL148 WL149 WL150 WL151 WL152 WL153 WL154 WL155 WL156 WL157 WL158 WL159 WL160 WL161 WL162
+ WL163 WL164 WL165 WL166 WL167 WL168 WL169 WL170 WL171 WL172 WL173 WL174 WL175 WL176 WL177 WL178 WL179
+ WL180 WL181 WL182 WL183 WL184 WL185 WL186 WL187 WL188 WL189 WL190 WL191 WL192 WL193 WL194 WL195 WL196
+ WL197 WL198 WL199 WL200 WL201 WL202 WL203 WL204 WL205 WL206 WL207 WL208 WL209 WL210 WL211 WL212 WL213
+ WL214 WL215 WL216 WL217 WL218 WL219 WL220 WL221 WL222 WL223 WL224 WL225 WL226 WL227 WL228 WL229 WL230
+ WL231 WL232 WL233 WL234 WL235 WL236 WL237 WL238 WL239 WL240 WL241 WL242 WL243 WL244 WL245 WL246 WL247
+ WL248 WL249 WL250 WL251 WL252 WL253 WL254 WL255 WL256 WL257 WL258 WL259 WL260 WL261 WL262 WL263 WL264
+ WL265 WL266 WL267 WL268 WL269 WL270 WL271 WL272 WL273 WL274 WL275 WL276 WL277 WL278 WL279 WL280 WL281
+ WL282 WL283 WL284 WL285 WL286 WL287 WL288 WL289 WL290 WL291 WL292 WL293 WL294 WL295 WL296 WL297 WL298
+ WL299 WL300 WL301 WL302 WL303 WL304 WL305 WL306 WL307 WL308 WL309 WL310 WL311 WL312 WL313 WL314 WL315
+ WL316 WL317 WL318 WL319 WL320 WL321 WL322 WL323 WL324 WL325 WL326 WL327 WL328 WL329 WL330 WL331 WL332
+ WL333 WL334 WL335 WL336 WL337 WL338 WL339 WL340 WL341 WL342 WL343 WL344 WL345 WL346 WL347 WL348 WL349
+ WL350 WL351 WL352 WL353 WL354 WL355 WL356 WL357 WL358 WL359 WL360 WL361 WL362 WL363 WL364 WL365 WL366
+ WL367 WL368 WL369 WL370 WL371 WL372 WL373 WL374 WL375 WL376 WL377 WL378 WL379 WL380 WL381 WL382 WL383
+ WL384 WL385 WL386 WL387 WL388 WL389 WL390 WL391 WL392 WL393 WL394 WL395 WL396 WL397 WL398 WL399 WL400
+ WL401 WL402 WL403 WL404 WL405 WL406 WL407 WL408 WL409 WL410 WL411 WL412 WL413 WL414 WL415 WL416 WL417
+ WL418 WL419 WL420 WL421 WL422 WL423 WL424 WL425 WL426 WL427 WL428 WL429 WL430 WL431 WL432 WL433 WL434
+ WL435 WL436 WL437 WL438 WL439 WL440 WL441 WL442 WL443 WL444 WL445 WL446 WL447 WL448 WL449 WL450 WL451
+ WL452 WL453 WL454 WL455 WL456 WL457 WL458 WL459 WL460 WL461 WL462 WL463 WL464 WL465 WL466 WL467 WL468
+ WL469 WL470 WL471 WL472 WL473 WL474 WL475 WL476 WL477 WL478 WL479 WL480 WL481 WL482 WL483 WL484 WL485
+ WL486 WL487 WL488 WL489 WL490 WL491 WL492 WL493 WL494 WL495 WL496 WL497 WL498 WL499 WL500 WL501 WL502
+ WL503 WL504 WL505 WL506 WL507 WL508 WL509 WL510 WL511 WL512 WL513 WL514 WL515 WL516 WL517 WL518 WL519
+ WL520 WL521 WL522 WL523 WL524 WL525 WL526 WL527 WL528 WL529 WL530 WL531 WL532 WL533 WL534 WL535 WL536
+ WL537 WL538 WL539 WL540 WL541 WL542 WL543 WL544 WL545 WL546 WL547 WL548 WL549 WL550 WL551 WL552 WL553
+ WL554 WL555 WL556 WL557 WL558 WL559 WL560 WL561 WL562 WL563 WL564 WL565 WL566 WL567 WL568 WL569 WL570
+ WL571 WL572 WL573 WL574 WL575 WL576 WL577 WL578 WL579 WL580 WL581 WL582 WL583 WL584 WL585 WL586 WL587
+ WL588 WL589 WL590 WL591 WL592 WL593 WL594 WL595 WL596 WL597 WL598 WL599 WL600 WL601 WL602 WL603 WL604
+ WL605 WL606 WL607 WL608 WL609 WL610 WL611 WL612 WL613 WL614 WL615 WL616 WL617 WL618 WL619 WL620 WL621
+ WL622 WL623 WL624 WL625 WL626 WL627 WL628 WL629 WL630 WL631 WL632 WL633 WL634 WL635 WL636 WL637 WL638
+ WL639 WL640 WL641 WL642 WL643 WL644 WL645 WL646 WL647 WL648 WL649 WL650 WL651 WL652 WL653 WL654 WL655
+ WL656 WL657 WL658 WL659 WL660 WL661 WL662 WL663 WL664 WL665 WL666 WL667 WL668 WL669 WL670 WL671 WL672
+ WL673 WL674 WL675 WL676 WL677 WL678 WL679 WL680 WL681 WL682 WL683 WL684 WL685 WL686 WL687 WL688 WL689
+ WL690 WL691 WL692 WL693 WL694 WL695 WL696 WL697 WL698 WL699 WL700 WL701 WL702 WL703 WL704 WL705 WL706
+ WL707 WL708 WL709 WL710 WL711 WL712 WL713 WL714 WL715 WL716 WL717 WL718 WL719 WL720 WL721 WL722 WL723
+ WL724 WL725 WL726 WL727 WL728 WL729 WL730 WL731 WL732 WL733 WL734 WL735 WL736 WL737 WL738 WL739 WL740
+ WL741 WL742 WL743 WL744 WL745 WL746 WL747 WL748 WL749 WL750 WL751 WL752 WL753 WL754 WL755 WL756 WL757
+ WL758 WL759 WL760 WL761 WL762 WL763 WL764 WL765 WL766 WL767 WL768 WL769 WL770 WL771 WL772 WL773 WL774
+ WL775 WL776 WL777 WL778 WL779 WL780 WL781 WL782 WL783 WL784 WL785 WL786 WL787 WL788 WL789 WL790 WL791
+ WL792 WL793 WL794 WL795 WL796 WL797 WL798 WL799 WL800 WL801 WL802 WL803 WL804 WL805 WL806 WL807 WL808
+ WL809 WL810 WL811 WL812 WL813 WL814 WL815 WL816 WL817 WL818 WL819 WL820 WL821 WL822 WL823 WL824 WL825
+ WL826 WL827 WL828 WL829 WL830 WL831 WL832 WL833 WL834 WL835 WL836 WL837 WL838 WL839 WL840 WL841 WL842
+ WL843 WL844 WL845 WL846 WL847 WL848 WL849 WL850 WL851 WL852 WL853 WL854 WL855 WL856 WL857 WL858 WL859
+ WL860 WL861 WL862 WL863 WL864 WL865 WL866 WL867 WL868 WL869 WL870 WL871 WL872 WL873 WL874 WL875 WL876
+ WL877 WL878 WL879 WL880 WL881 WL882 WL883 WL884 WL885 WL886 WL887 WL888 WL889 WL890 WL891 WL892 WL893
+ WL894 WL895 WL896 WL897 WL898 WL899 WL900 WL901 WL902 WL903 WL904 WL905 WL906 WL907 WL908 WL909 WL910
+ WL911 WL912 WL913 WL914 WL915 WL916 WL917 WL918 WL919 WL920 WL921 WL922 WL923 WL924 WL925 WL926 WL927
+ WL928 WL929 WL930 WL931 WL932 WL933 WL934 WL935 WL936 WL937 WL938 WL939 WL940 WL941 WL942 WL943 WL944
+ WL945 WL946 WL947 WL948 WL949 WL950 WL951 WL952 WL953 WL954 WL955 WL956 WL957 WL958 WL959 WL960 WL961
+ WL962 WL963 WL964 WL965 WL966 WL967 WL968 WL969 WL970 WL971 WL972 WL973 WL974 WL975 WL976 WL977 WL978
+ WL979 WL980 WL981 WL982 WL983 WL984 WL985 WL986 WL987 WL988 WL989 WL990 WL991 WL992 WL993 WL994 WL995
+ WL996 WL997 WL998 WL999 WL1000 WL1001 WL1002 WL1003 WL1004 WL1005 WL1006 WL1007 WL1008 WL1009 WL1010
+ WL1011 WL1012 WL1013 WL1014 WL1015 WL1016 WL1017 WL1018 WL1019 WL1020 WL1021 WL1022 WL1023
+ 32x1024_truncation_sram
x2 net63 Read31 net61 Read30 Read29 net59 Read28 net57 net55 Read27 Read26 net35 Read25 net33 net54
+ Read24 net64 net62 net60 Trunk31 net58 Trunk30 net56 net37 Trunk29 Trunk28 net36 net34 Trunk27 Trunk26
+ DataOut31 Trunk25 DataOut30 Trunk24 DataOut29 DataOut28 DataOut27 DataOut26 DataOut25 Byte_Mode_EnableBar
+ DataOut24 tail_IO3 Tail_In vssd1 vccd1 1bytetruncationmanagerwithand
x3 net32 Read23 net30 Read22 Read21 net28 Read20 net26 net24 Read19 Read18 net22 Read17 net20 net18
+ Read16 net31 net29 net27 Trunk23 net25 Trunk22 net23 net21 Trunk21 Trunk20 net19 net17 Trunk19 Trunk18
+ DataOut23 Trunk17 DataOut22 Trunk16 DataOut21 DataOut20 DataOut19 DataOut18 DataOut17 Byte_Mode_EnableBar
+ DataOut16 tail_IO2 tail_IO3 vssd1 vccd1 1bytetruncationmanagerwithand
x4 net16 Read15 net14 Read14 Read13 net12 Read12 net10 net8 Read11 Read10 net6 Read9 net4 net2 Read8
+ net15 net13 net11 Trunk15 net9 Trunk14 net7 net5 Trunk13 Trunk12 net3 net1 Trunk11 Trunk10 DataOut15
+ Trunk9 DataOut14 Trunk8 DataOut13 DataOut12 DataOut11 DataOut10 DataOut9 Byte_Mode_EnableBar DataOut8
+ tail_IO1 tail_IO2 vssd1 vccd1 1bytetruncationmanagerwithand
x5 net52 Read7 net50 Read6 Read5 net48 Read4 net46 net44 Read3 Read2 net42 Read1 net40 net38 Read0
+ net53 net51 net49 Trunk7 net47 Trunk6 net45 net43 Trunk5 Trunk4 net41 net39 Trunk3 Trunk2 DataOut7 Trunk1
+ DataOut6 Trunk0 DataOut5 DataOut4 DataOut3 DataOut2 DataOut1 Byte_Mode_EnableBar DataOut0 Tail_Out tail_IO1
+ vssd1 vccd1 1bytetruncationmanagerwithand
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/32x1024_truncation_sram.sym
*+ # of pins=1157
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/32x1024_truncation_sram.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/32x1024_truncation_sram.sch
.subckt 32x1024_truncation_sram vcc vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3
+ vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10
+ gnd_bl10 vcc_bl11 gnd_bl11 vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16
+ gnd_bl16 vcc_bl17 gnd_bl17 vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22
+ gnd_bl22 vcc_bl23 gnd_bl23 vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28
+ gnd_bl28 vcc_bl29 gnd_bl29 vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 gnd PRE writeen readen DataIn31 DataIn30
+ DataIn29 DataIn28 DataIn27 DataIn26 DataIn25 DataIn24 DataIn23 DataIn22 DataIn21 DataIn20 DataIn19 DataIn18
+ DataIn17 DataIn16 DataIn15 DataIn14 DataIn13 DataIn12 DataIn11 DataIn10 DataIn9 DataIn8 DataIn7 DataIn6
+ DataIn5 DataIn4 DataIn3 DataIn2 DataIn1 DataIn0 DataOut31 DataOut30 DataOut29 DataOut28 DataOut27 DataOut26
+ DataOut25 DataOut24 DataOut23 DataOut22 DataOut21 DataOut20 DataOut19 DataOut18 DataOut17 DataOut16 DataOut15
+ DataOut14 DataOut13 DataOut12 DataOut11 DataOut10 DataOut9 DataOut8 DataOut7 DataOut6 DataOut5 DataOut4
+ DataOut3 DataOut2 DataOut1 DataOut0 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15
+ WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36
+ WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57
+ WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78
+ WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99
+ WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116
+ WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 WL128 WL129 WL130 WL131 WL132 WL133
+ WL134 WL135 WL136 WL137 WL138 WL139 WL140 WL141 WL142 WL143 WL144 WL145 WL146 WL147 WL148 WL149 WL150
+ WL151 WL152 WL153 WL154 WL155 WL156 WL157 WL158 WL159 WL160 WL161 WL162 WL163 WL164 WL165 WL166 WL167
+ WL168 WL169 WL170 WL171 WL172 WL173 WL174 WL175 WL176 WL177 WL178 WL179 WL180 WL181 WL182 WL183 WL184
+ WL185 WL186 WL187 WL188 WL189 WL190 WL191 WL192 WL193 WL194 WL195 WL196 WL197 WL198 WL199 WL200 WL201
+ WL202 WL203 WL204 WL205 WL206 WL207 WL208 WL209 WL210 WL211 WL212 WL213 WL214 WL215 WL216 WL217 WL218
+ WL219 WL220 WL221 WL222 WL223 WL224 WL225 WL226 WL227 WL228 WL229 WL230 WL231 WL232 WL233 WL234 WL235
+ WL236 WL237 WL238 WL239 WL240 WL241 WL242 WL243 WL244 WL245 WL246 WL247 WL248 WL249 WL250 WL251 WL252
+ WL253 WL254 WL255 WL256 WL257 WL258 WL259 WL260 WL261 WL262 WL263 WL264 WL265 WL266 WL267 WL268 WL269
+ WL270 WL271 WL272 WL273 WL274 WL275 WL276 WL277 WL278 WL279 WL280 WL281 WL282 WL283 WL284 WL285 WL286
+ WL287 WL288 WL289 WL290 WL291 WL292 WL293 WL294 WL295 WL296 WL297 WL298 WL299 WL300 WL301 WL302 WL303
+ WL304 WL305 WL306 WL307 WL308 WL309 WL310 WL311 WL312 WL313 WL314 WL315 WL316 WL317 WL318 WL319 WL320
+ WL321 WL322 WL323 WL324 WL325 WL326 WL327 WL328 WL329 WL330 WL331 WL332 WL333 WL334 WL335 WL336 WL337
+ WL338 WL339 WL340 WL341 WL342 WL343 WL344 WL345 WL346 WL347 WL348 WL349 WL350 WL351 WL352 WL353 WL354
+ WL355 WL356 WL357 WL358 WL359 WL360 WL361 WL362 WL363 WL364 WL365 WL366 WL367 WL368 WL369 WL370 WL371
+ WL372 WL373 WL374 WL375 WL376 WL377 WL378 WL379 WL380 WL381 WL382 WL383 WL384 WL385 WL386 WL387 WL388
+ WL389 WL390 WL391 WL392 WL393 WL394 WL395 WL396 WL397 WL398 WL399 WL400 WL401 WL402 WL403 WL404 WL405
+ WL406 WL407 WL408 WL409 WL410 WL411 WL412 WL413 WL414 WL415 WL416 WL417 WL418 WL419 WL420 WL421 WL422
+ WL423 WL424 WL425 WL426 WL427 WL428 WL429 WL430 WL431 WL432 WL433 WL434 WL435 WL436 WL437 WL438 WL439
+ WL440 WL441 WL442 WL443 WL444 WL445 WL446 WL447 WL448 WL449 WL450 WL451 WL452 WL453 WL454 WL455 WL456
+ WL457 WL458 WL459 WL460 WL461 WL462 WL463 WL464 WL465 WL466 WL467 WL468 WL469 WL470 WL471 WL472 WL473
+ WL474 WL475 WL476 WL477 WL478 WL479 WL480 WL481 WL482 WL483 WL484 WL485 WL486 WL487 WL488 WL489 WL490
+ WL491 WL492 WL493 WL494 WL495 WL496 WL497 WL498 WL499 WL500 WL501 WL502 WL503 WL504 WL505 WL506 WL507
+ WL508 WL509 WL510 WL511 WL512 WL513 WL514 WL515 WL516 WL517 WL518 WL519 WL520 WL521 WL522 WL523 WL524
+ WL525 WL526 WL527 WL528 WL529 WL530 WL531 WL532 WL533 WL534 WL535 WL536 WL537 WL538 WL539 WL540 WL541
+ WL542 WL543 WL544 WL545 WL546 WL547 WL548 WL549 WL550 WL551 WL552 WL553 WL554 WL555 WL556 WL557 WL558
+ WL559 WL560 WL561 WL562 WL563 WL564 WL565 WL566 WL567 WL568 WL569 WL570 WL571 WL572 WL573 WL574 WL575
+ WL576 WL577 WL578 WL579 WL580 WL581 WL582 WL583 WL584 WL585 WL586 WL587 WL588 WL589 WL590 WL591 WL592
+ WL593 WL594 WL595 WL596 WL597 WL598 WL599 WL600 WL601 WL602 WL603 WL604 WL605 WL606 WL607 WL608 WL609
+ WL610 WL611 WL612 WL613 WL614 WL615 WL616 WL617 WL618 WL619 WL620 WL621 WL622 WL623 WL624 WL625 WL626
+ WL627 WL628 WL629 WL630 WL631 WL632 WL633 WL634 WL635 WL636 WL637 WL638 WL639 WL640 WL641 WL642 WL643
+ WL644 WL645 WL646 WL647 WL648 WL649 WL650 WL651 WL652 WL653 WL654 WL655 WL656 WL657 WL658 WL659 WL660
+ WL661 WL662 WL663 WL664 WL665 WL666 WL667 WL668 WL669 WL670 WL671 WL672 WL673 WL674 WL675 WL676 WL677
+ WL678 WL679 WL680 WL681 WL682 WL683 WL684 WL685 WL686 WL687 WL688 WL689 WL690 WL691 WL692 WL693 WL694
+ WL695 WL696 WL697 WL698 WL699 WL700 WL701 WL702 WL703 WL704 WL705 WL706 WL707 WL708 WL709 WL710 WL711
+ WL712 WL713 WL714 WL715 WL716 WL717 WL718 WL719 WL720 WL721 WL722 WL723 WL724 WL725 WL726 WL727 WL728
+ WL729 WL730 WL731 WL732 WL733 WL734 WL735 WL736 WL737 WL738 WL739 WL740 WL741 WL742 WL743 WL744 WL745
+ WL746 WL747 WL748 WL749 WL750 WL751 WL752 WL753 WL754 WL755 WL756 WL757 WL758 WL759 WL760 WL761 WL762
+ WL763 WL764 WL765 WL766 WL767 WL768 WL769 WL770 WL771 WL772 WL773 WL774 WL775 WL776 WL777 WL778 WL779
+ WL780 WL781 WL782 WL783 WL784 WL785 WL786 WL787 WL788 WL789 WL790 WL791 WL792 WL793 WL794 WL795 WL796
+ WL797 WL798 WL799 WL800 WL801 WL802 WL803 WL804 WL805 WL806 WL807 WL808 WL809 WL810 WL811 WL812 WL813
+ WL814 WL815 WL816 WL817 WL818 WL819 WL820 WL821 WL822 WL823 WL824 WL825 WL826 WL827 WL828 WL829 WL830
+ WL831 WL832 WL833 WL834 WL835 WL836 WL837 WL838 WL839 WL840 WL841 WL842 WL843 WL844 WL845 WL846 WL847
+ WL848 WL849 WL850 WL851 WL852 WL853 WL854 WL855 WL856 WL857 WL858 WL859 WL860 WL861 WL862 WL863 WL864
+ WL865 WL866 WL867 WL868 WL869 WL870 WL871 WL872 WL873 WL874 WL875 WL876 WL877 WL878 WL879 WL880 WL881
+ WL882 WL883 WL884 WL885 WL886 WL887 WL888 WL889 WL890 WL891 WL892 WL893 WL894 WL895 WL896 WL897 WL898
+ WL899 WL900 WL901 WL902 WL903 WL904 WL905 WL906 WL907 WL908 WL909 WL910 WL911 WL912 WL913 WL914 WL915
+ WL916 WL917 WL918 WL919 WL920 WL921 WL922 WL923 WL924 WL925 WL926 WL927 WL928 WL929 WL930 WL931 WL932
+ WL933 WL934 WL935 WL936 WL937 WL938 WL939 WL940 WL941 WL942 WL943 WL944 WL945 WL946 WL947 WL948 WL949
+ WL950 WL951 WL952 WL953 WL954 WL955 WL956 WL957 WL958 WL959 WL960 WL961 WL962 WL963 WL964 WL965 WL966
+ WL967 WL968 WL969 WL970 WL971 WL972 WL973 WL974 WL975 WL976 WL977 WL978 WL979 WL980 WL981 WL982 WL983
+ WL984 WL985 WL986 WL987 WL988 WL989 WL990 WL991 WL992 WL993 WL994 WL995 WL996 WL997 WL998 WL999 WL1000
+ WL1001 WL1002 WL1003 WL1004 WL1005 WL1006 WL1007 WL1008 WL1009 WL1010 WL1011 WL1012 WL1013 WL1014 WL1015
+ WL1016 WL1017 WL1018 WL1019 WL1020 WL1021 WL1022 WL1023
*.PININFO vcc_bl0:B vcc_bl1:B vcc_bl2:B vcc_bl3:B gnd_bl0:B gnd_bl1:B gnd_bl2:B gnd_bl3:B vcc_bl4:B
*+ vcc_bl5:B vcc_bl6:B vcc_bl7:B gnd_bl4:B gnd_bl5:B gnd_bl6:B gnd_bl7:B vcc_bl8:B vcc_bl9:B vcc_bl10:B
*+ vcc_bl11:B gnd_bl8:B gnd_bl9:B gnd_bl10:B gnd_bl11:B vcc_bl12:B vcc_bl13:B vcc_bl14:B vcc_bl15:B gnd_bl12:B
*+ gnd_bl13:B gnd_bl14:B gnd_bl15:B vcc_bl16:B vcc_bl17:B vcc_bl18:B vcc_bl19:B gnd_bl16:B gnd_bl17:B gnd_bl18:B
*+ gnd_bl19:B vcc_bl20:B vcc_bl21:B vcc_bl22:B vcc_bl23:B gnd_bl20:B gnd_bl21:B gnd_bl22:B gnd_bl23:B vcc_bl24:B
*+ vcc_bl25:B vcc_bl26:B vcc_bl27:B gnd_bl24:B gnd_bl25:B gnd_bl26:B gnd_bl27:B vcc_bl28:B vcc_bl29:B vcc_bl30:B
*+ vcc_bl31:B gnd_bl28:B gnd_bl29:B gnd_bl30:B gnd_bl31:B gnd:B WL160:I WL161:I WL162:I WL163:I WL164:I WL165:I
*+ WL166:I WL167:I WL168:I WL169:I WL170:I WL171:I WL172:I WL173:I WL174:I WL175:I WL176:I WL177:I WL178:I
*+ WL179:I WL180:I WL181:I WL182:I WL183:I WL184:I WL185:I WL186:I WL187:I WL188:I WL189:I WL190:I WL191:I
*+ WL224:I WL225:I WL226:I WL227:I WL228:I WL229:I WL230:I WL231:I WL232:I WL233:I WL234:I WL235:I WL236:I
*+ WL237:I WL238:I WL239:I WL240:I WL241:I WL242:I WL243:I WL244:I WL245:I WL246:I WL247:I WL248:I WL249:I
*+ WL250:I WL251:I WL252:I WL253:I WL254:I WL255:I WL256:I WL257:I WL258:I WL259:I WL260:I WL261:I WL262:I
*+ WL263:I WL264:I WL265:I WL266:I WL267:I WL268:I WL269:I WL270:I WL271:I WL272:I WL273:I WL274:I WL275:I
*+ WL276:I WL277:I WL278:I WL279:I WL280:I WL281:I WL282:I WL283:I WL284:I WL285:I WL286:I WL287:I WL288:I
*+ WL289:I WL290:I WL291:I WL292:I WL293:I WL294:I WL295:I WL296:I WL297:I WL298:I WL299:I WL300:I WL301:I
*+ WL302:I WL303:I WL304:I WL305:I WL306:I WL307:I WL308:I WL309:I WL310:I WL311:I WL312:I WL313:I WL314:I
*+ WL315:I WL316:I WL317:I WL318:I WL319:I WL320:I WL321:I WL322:I WL323:I WL324:I WL325:I WL326:I WL327:I
*+ WL328:I WL329:I WL330:I WL331:I WL332:I WL333:I WL334:I WL335:I WL336:I WL337:I WL338:I WL339:I WL340:I
*+ WL341:I WL342:I WL343:I WL344:I WL345:I WL346:I WL347:I WL348:I WL349:I WL350:I WL351:I WL352:I WL353:I
*+ WL354:I WL355:I WL356:I WL357:I WL358:I WL359:I WL360:I WL361:I WL362:I WL363:I WL364:I WL365:I WL366:I
*+ WL367:I WL368:I WL369:I WL370:I WL371:I WL372:I WL373:I WL374:I WL375:I WL376:I WL377:I WL378:I WL379:I
*+ WL380:I WL381:I WL382:I WL383:I WL384:I WL385:I WL386:I WL387:I WL388:I WL389:I WL390:I WL391:I WL392:I
*+ WL393:I WL394:I WL395:I WL396:I WL397:I WL398:I WL399:I WL400:I WL401:I WL402:I WL403:I WL404:I WL405:I
*+ WL406:I WL407:I WL408:I WL409:I WL410:I WL411:I WL412:I WL413:I WL414:I WL415:I WL416:I WL417:I WL418:I
*+ WL419:I WL420:I WL421:I WL422:I WL423:I WL424:I WL425:I WL426:I WL427:I WL428:I WL429:I WL430:I WL431:I
*+ WL432:I WL433:I WL434:I WL435:I WL436:I WL437:I WL438:I WL439:I WL440:I WL441:I WL442:I WL443:I WL444:I
*+ WL445:I WL446:I WL447:I WL448:I WL449:I WL450:I WL451:I WL452:I WL453:I WL454:I WL455:I WL456:I WL457:I
*+ WL458:I WL459:I WL460:I WL461:I WL462:I WL463:I WL464:I WL465:I WL466:I WL467:I WL468:I WL469:I WL470:I
*+ WL471:I WL472:I WL473:I WL474:I WL475:I WL476:I WL477:I WL478:I WL479:I WL480:I WL481:I WL482:I WL483:I
*+ WL484:I WL485:I WL486:I WL487:I WL488:I WL489:I WL490:I WL491:I WL492:I WL493:I WL494:I WL495:I WL496:I
*+ WL497:I WL498:I WL499:I WL500:I WL501:I WL502:I WL503:I WL504:I WL505:I WL506:I WL507:I WL508:I WL509:I
*+ WL510:I WL511:I WL512:I WL513:I WL514:I WL515:I WL516:I WL517:I WL518:I WL519:I WL520:I WL521:I WL522:I
*+ WL523:I WL524:I WL525:I WL526:I WL527:I WL528:I WL529:I WL530:I WL531:I WL532:I WL533:I WL534:I WL535:I
*+ WL536:I WL537:I WL538:I WL539:I WL540:I WL541:I WL542:I WL543:I WL544:I WL545:I WL546:I WL547:I WL548:I
*+ WL549:I WL550:I WL551:I WL552:I WL553:I WL554:I WL555:I WL556:I WL557:I WL558:I WL559:I WL560:I WL561:I
*+ WL562:I WL563:I WL564:I WL565:I WL566:I WL567:I WL568:I WL569:I WL570:I WL571:I WL572:I WL573:I WL574:I
*+ WL575:I WL576:I WL577:I WL578:I WL579:I WL580:I WL581:I WL582:I WL583:I WL584:I WL585:I WL586:I WL587:I
*+ WL588:I WL589:I WL590:I WL591:I WL592:I WL593:I WL594:I WL595:I WL596:I WL597:I WL598:I WL599:I WL600:I
*+ WL601:I WL602:I WL603:I WL604:I WL605:I WL606:I WL607:I WL608:I WL609:I WL610:I WL611:I WL612:I WL613:I
*+ WL614:I WL615:I WL616:I WL617:I WL618:I WL619:I WL620:I WL621:I WL622:I WL623:I WL624:I WL625:I WL626:I
*+ WL627:I WL628:I WL629:I WL630:I WL631:I WL632:I WL633:I WL634:I WL635:I WL636:I WL637:I WL638:I WL639:I
*+ WL640:I WL641:I WL642:I WL643:I WL644:I WL645:I WL646:I WL647:I WL648:I WL649:I WL650:I WL651:I WL652:I
*+ WL653:I WL654:I WL655:I WL656:I WL657:I WL658:I WL659:I WL660:I WL661:I WL662:I WL663:I WL664:I WL665:I
*+ WL666:I WL667:I WL668:I WL669:I WL670:I WL671:I WL672:I WL673:I WL674:I WL675:I WL676:I WL677:I WL678:I
*+ WL679:I WL680:I WL681:I WL682:I WL683:I WL684:I WL685:I WL686:I WL687:I WL688:I WL689:I WL690:I WL691:I
*+ WL692:I WL693:I WL694:I WL695:I WL696:I WL697:I WL698:I WL699:I WL700:I WL701:I WL702:I WL703:I WL704:I
*+ WL705:I WL706:I WL707:I WL708:I WL709:I WL710:I WL711:I WL712:I WL713:I WL714:I WL715:I WL716:I WL717:I
*+ WL718:I WL719:I WL720:I WL721:I WL722:I WL723:I WL724:I WL725:I WL726:I WL727:I WL728:I WL729:I WL730:I
*+ WL731:I WL732:I WL733:I WL734:I WL735:I WL736:I WL737:I WL738:I WL739:I WL740:I WL741:I WL742:I WL743:I
*+ WL744:I WL745:I WL746:I WL747:I WL748:I WL749:I WL750:I WL751:I WL752:I WL753:I WL754:I WL755:I WL756:I
*+ WL757:I WL758:I WL759:I WL760:I WL761:I WL762:I WL763:I WL764:I WL765:I WL766:I WL767:I WL768:I WL769:I
*+ WL770:I WL771:I WL772:I WL773:I WL774:I WL775:I WL776:I WL777:I WL778:I WL779:I WL780:I WL781:I WL782:I
*+ WL783:I WL784:I WL785:I WL786:I WL787:I WL788:I WL789:I WL790:I WL791:I WL792:I WL793:I WL794:I WL795:I
*+ WL796:I WL797:I WL798:I WL799:I WL800:I WL801:I WL802:I WL803:I WL804:I WL805:I WL806:I WL807:I WL808:I
*+ WL809:I WL810:I WL811:I WL812:I WL813:I WL814:I WL815:I WL816:I WL817:I WL818:I WL819:I WL820:I WL821:I
*+ WL822:I WL823:I WL824:I WL825:I WL826:I WL827:I WL828:I WL829:I WL830:I WL831:I WL832:I WL833:I WL834:I
*+ WL835:I WL836:I WL837:I WL838:I WL839:I WL840:I WL841:I WL842:I WL843:I WL844:I WL845:I WL846:I WL847:I
*+ WL848:I WL849:I WL850:I WL851:I WL852:I WL853:I WL854:I WL855:I WL856:I WL857:I WL858:I WL859:I WL860:I
*+ WL861:I WL862:I WL863:I WL864:I WL865:I WL866:I WL867:I WL868:I WL869:I WL870:I WL871:I WL872:I WL873:I
*+ WL874:I WL875:I WL876:I WL877:I WL878:I WL879:I WL880:I WL881:I WL882:I WL883:I WL884:I WL885:I WL886:I
*+ WL887:I WL888:I WL889:I WL890:I WL891:I WL892:I WL893:I WL894:I WL895:I WL896:I WL897:I WL898:I WL899:I
*+ WL900:I WL901:I WL902:I WL903:I WL904:I WL905:I WL906:I WL907:I WL908:I WL909:I WL910:I WL911:I WL912:I
*+ WL913:I WL914:I WL915:I WL916:I WL917:I WL918:I WL919:I WL920:I WL921:I WL922:I WL923:I WL924:I WL925:I
*+ WL926:I WL927:I WL928:I WL929:I WL930:I WL931:I WL932:I WL933:I WL934:I WL935:I WL936:I WL937:I WL938:I
*+ WL939:I WL940:I WL941:I WL942:I WL943:I WL944:I WL945:I WL946:I WL947:I WL948:I WL949:I WL950:I WL951:I
*+ WL952:I WL953:I WL954:I WL955:I WL956:I WL957:I WL958:I WL959:I WL960:I WL961:I WL962:I WL963:I WL964:I
*+ WL965:I WL966:I WL967:I WL968:I WL969:I WL970:I WL971:I WL972:I WL973:I WL974:I WL975:I WL976:I WL977:I
*+ WL978:I WL979:I WL980:I WL981:I WL982:I WL983:I WL984:I WL985:I WL986:I WL987:I WL988:I WL989:I WL990:I
*+ WL991:I WL992:I WL993:I WL994:I WL995:I WL996:I WL997:I WL998:I WL999:I WL1000:I WL1001:I WL1002:I WL1003:I
*+ WL1004:I WL1005:I WL1006:I WL1007:I WL1008:I WL1009:I WL1010:I WL1011:I WL1012:I WL1013:I WL1014:I WL1015:I
*+ WL1016:I WL1017:I WL1018:I WL1019:I WL1020:I WL1021:I WL1022:I WL1023:I WL32:I WL33:I WL34:I WL35:I WL36:I
*+ WL37:I WL38:I WL39:I WL40:I WL41:I WL42:I WL43:I WL44:I WL45:I WL46:I WL47:I WL48:I WL49:I WL50:I WL51:I
*+ WL52:I WL53:I WL54:I WL55:I WL56:I WL57:I WL58:I WL59:I WL60:I WL61:I WL62:I WL63:I WL64:I WL65:I WL66:I
*+ WL67:I WL68:I WL69:I WL70:I WL71:I WL72:I WL73:I WL74:I WL75:I WL76:I WL77:I WL78:I WL79:I WL80:I WL81:I
*+ WL82:I WL83:I WL84:I WL85:I WL86:I WL87:I WL88:I WL89:I WL90:I WL91:I WL92:I WL93:I WL94:I WL95:I WL96:I
*+ WL97:I WL98:I WL99:I WL100:I WL101:I WL102:I WL103:I WL104:I WL105:I WL106:I WL107:I WL108:I WL109:I
*+ WL110:I WL111:I WL112:I WL113:I WL114:I WL115:I WL116:I WL117:I WL118:I WL119:I WL120:I WL121:I WL122:I
*+ WL123:I WL124:I WL125:I WL126:I WL127:I WL128:I WL129:I WL130:I WL131:I WL132:I WL133:I WL134:I WL135:I
*+ WL136:I WL137:I WL138:I WL139:I WL140:I WL141:I WL142:I WL143:I WL144:I WL145:I WL146:I WL147:I WL148:I
*+ WL149:I WL150:I WL151:I WL152:I WL153:I WL154:I WL155:I WL156:I WL157:I WL158:I WL159:I WL0:I WL1:I WL2:I
*+ WL3:I WL4:I WL5:I WL6:I WL7:I WL8:I WL9:I WL10:I WL11:I WL12:I WL13:I WL14:I WL15:I WL16:I WL17:I WL18:I
*+ WL19:I WL20:I WL21:I WL22:I WL23:I WL24:I WL25:I WL26:I WL27:I WL28:I WL29:I WL30:I WL31:I WL192:I WL193:I
*+ WL194:I WL195:I WL196:I WL197:I WL198:I WL199:I WL200:I WL201:I WL202:I WL203:I WL204:I WL205:I WL206:I
*+ WL207:I WL208:I WL209:I WL210:I WL211:I WL212:I WL213:I WL214:I WL215:I WL216:I WL217:I WL218:I WL219:I
*+ WL220:I WL221:I WL222:I WL223:I vcc:B PRE:I writeen:I readen:I DataIn30:I DataIn29:I DataIn28:I DataIn27:I
*+ DataIn26:I DataIn25:I DataIn24:I DataIn23:I DataIn22:I DataIn21:I DataIn20:I DataIn19:I DataIn18:I DataIn17:I
*+ DataIn16:I DataIn15:I DataIn14:I DataIn13:I DataIn12:I DataIn11:I DataIn10:I DataIn9:I DataIn8:I DataIn7:I
*+ DataIn6:I DataIn5:I DataIn4:I DataIn3:I DataIn2:I DataIn1:I DataIn0:I DataIn31:I DataOut30:O DataOut29:O
*+ DataOut28:O DataOut27:O DataOut26:O DataOut25:O DataOut24:O DataOut23:O DataOut22:O DataOut21:O DataOut20:O
*+ DataOut19:O DataOut18:O DataOut17:O DataOut16:O DataOut15:O DataOut14:O DataOut13:O DataOut12:O DataOut11:O
*+ DataOut10:O DataOut9:O DataOut8:O DataOut7:O DataOut6:O DataOut5:O DataOut4:O DataOut3:O DataOut2:O DataOut1:O
*+ DataOut0:O DataOut31:O
x98 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net1 net2 net3 net4 net5 net6 net7 net8 net9 net10 net11 net12 net13
+ net14 net15 net16 net17 net18 net19 net20 net21 net22 net23 net24 net25 net26 net27 net28 net29 net30
+ net31 net32 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31 Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28
+ Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23 Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20
+ Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25 Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29
+ Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x102 gnd WL32 net1 vcc buffer
x130 gnd WL33 net2 vcc buffer
x131 gnd WL34 net3 vcc buffer
x132 gnd WL35 net4 vcc buffer
x134 gnd WL36 net5 vcc buffer
x135 gnd WL37 net6 vcc buffer
x136 gnd WL38 net7 vcc buffer
x137 gnd WL39 net8 vcc buffer
x138 gnd WL40 net9 vcc buffer
x139 gnd WL41 net10 vcc buffer
x140 gnd WL42 net11 vcc buffer
x141 gnd WL43 net12 vcc buffer
x142 gnd WL44 net13 vcc buffer
x143 gnd WL45 net14 vcc buffer
x144 gnd WL46 net15 vcc buffer
x145 gnd WL47 net16 vcc buffer
x146 gnd WL48 net17 vcc buffer
x147 gnd WL49 net18 vcc buffer
x148 gnd WL50 net19 vcc buffer
x149 gnd WL51 net20 vcc buffer
x150 gnd WL52 net21 vcc buffer
x151 gnd WL53 net22 vcc buffer
x152 gnd WL54 net23 vcc buffer
x153 gnd WL55 net24 vcc buffer
x154 gnd WL56 net25 vcc buffer
x155 gnd WL57 net26 vcc buffer
x156 gnd WL58 net27 vcc buffer
x157 gnd WL59 net28 vcc buffer
x158 gnd WL60 net29 vcc buffer
x159 gnd WL61 net30 vcc buffer
x160 gnd WL62 net31 vcc buffer
x161 gnd WL63 net32 vcc buffer
x5 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net33 net34 net35 net36 net37 net38 net39 net40 net41 net42 net43 net44
+ net45 net46 net47 net48 net49 net50 net51 net52 net53 net54 net55 net56 net57 net58 net59 net60 net61
+ net62 net63 net64 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31 Bl31 Blb30 Blb7 Bl7 Blb6 Bl6
+ Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23 Blb22 Bl3 Blb2 Blb21 Blb20 Bl2
+ Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25 Bl26 Bl16 Bl27 Blb15 Bl28 Bl15
+ Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x103 gnd WL0 net33 vcc buffer
x104 gnd WL1 net34 vcc buffer
x105 gnd WL2 net35 vcc buffer
x106 gnd WL3 net36 vcc buffer
x107 gnd WL4 net37 vcc buffer
x108 gnd WL5 net38 vcc buffer
x109 gnd WL6 net39 vcc buffer
x110 gnd WL7 net40 vcc buffer
x111 gnd WL8 net41 vcc buffer
x112 gnd WL9 net42 vcc buffer
x113 gnd WL10 net43 vcc buffer
x114 gnd WL11 net44 vcc buffer
x115 gnd WL12 net45 vcc buffer
x116 gnd WL13 net46 vcc buffer
x117 gnd WL14 net47 vcc buffer
x118 gnd WL15 net48 vcc buffer
x119 gnd WL16 net49 vcc buffer
x120 gnd WL17 net50 vcc buffer
x121 gnd WL18 net51 vcc buffer
x122 gnd WL19 net52 vcc buffer
x123 gnd WL20 net53 vcc buffer
x124 gnd WL21 net54 vcc buffer
x125 gnd WL22 net55 vcc buffer
x126 gnd WL23 net56 vcc buffer
x127 gnd WL24 net57 vcc buffer
x128 gnd WL25 net58 vcc buffer
x129 gnd WL26 net59 vcc buffer
x193 gnd WL27 net60 vcc buffer
x194 gnd WL28 net61 vcc buffer
x195 gnd WL29 net62 vcc buffer
x196 gnd WL30 net63 vcc buffer
x197 gnd WL31 net64 vcc buffer
x99 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net65 net66 net67 net68 net69 net70 net71 net72 net73 net74 net75 net76
+ net77 net78 net79 net80 net81 net82 net83 net84 net85 net86 net87 net88 net89 net90 net91 net92 net93
+ net94 net95 net96 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31 Bl31 Blb30 Blb7 Bl7 Blb6 Bl6
+ Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23 Blb22 Bl3 Blb2 Blb21 Blb20 Bl2
+ Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25 Bl26 Bl16 Bl27 Blb15 Bl28 Bl15
+ Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x100 gnd WL64 net65 vcc buffer
x101 gnd WL65 net66 vcc buffer
x133 gnd WL66 net67 vcc buffer
x162 gnd WL67 net68 vcc buffer
x163 gnd WL68 net69 vcc buffer
x164 gnd WL69 net70 vcc buffer
x165 gnd WL70 net71 vcc buffer
x166 gnd WL71 net72 vcc buffer
x167 gnd WL72 net73 vcc buffer
x168 gnd WL73 net74 vcc buffer
x169 gnd WL74 net75 vcc buffer
x170 gnd WL75 net76 vcc buffer
x171 gnd WL76 net77 vcc buffer
x172 gnd WL77 net78 vcc buffer
x173 gnd WL78 net79 vcc buffer
x174 gnd WL79 net80 vcc buffer
x175 gnd WL80 net81 vcc buffer
x176 gnd WL81 net82 vcc buffer
x177 gnd WL82 net83 vcc buffer
x178 gnd WL83 net84 vcc buffer
x179 gnd WL84 net85 vcc buffer
x180 gnd WL85 net86 vcc buffer
x181 gnd WL86 net87 vcc buffer
x182 gnd WL87 net88 vcc buffer
x183 gnd WL88 net89 vcc buffer
x184 gnd WL89 net90 vcc buffer
x185 gnd WL90 net91 vcc buffer
x186 gnd WL91 net92 vcc buffer
x187 gnd WL92 net93 vcc buffer
x188 gnd WL93 net94 vcc buffer
x189 gnd WL94 net95 vcc buffer
x190 gnd WL95 net96 vcc buffer
x191 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net97 net98 net99 net100 net101 net102 net103 net104 net105 net106
+ net107 net108 net109 net110 net111 net112 net113 net114 net115 net116 net117 net118 net119 net120 net121
+ net122 net123 net124 net125 net126 net127 net128 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x192 gnd WL96 net97 vcc buffer
x198 gnd WL97 net98 vcc buffer
x199 gnd WL98 net99 vcc buffer
x200 gnd WL99 net100 vcc buffer
x201 gnd WL100 net101 vcc buffer
x202 gnd WL101 net102 vcc buffer
x203 gnd WL102 net103 vcc buffer
x204 gnd WL103 net104 vcc buffer
x205 gnd WL104 net105 vcc buffer
x206 gnd WL105 net106 vcc buffer
x207 gnd WL106 net107 vcc buffer
x208 gnd WL107 net108 vcc buffer
x209 gnd WL108 net109 vcc buffer
x210 gnd WL109 net110 vcc buffer
x211 gnd WL110 net111 vcc buffer
x212 gnd WL111 net112 vcc buffer
x213 gnd WL112 net113 vcc buffer
x214 gnd WL113 net114 vcc buffer
x215 gnd WL114 net115 vcc buffer
x216 gnd WL115 net116 vcc buffer
x217 gnd WL116 net117 vcc buffer
x218 gnd WL117 net118 vcc buffer
x219 gnd WL118 net119 vcc buffer
x220 gnd WL119 net120 vcc buffer
x221 gnd WL120 net121 vcc buffer
x222 gnd WL121 net122 vcc buffer
x223 gnd WL122 net123 vcc buffer
x224 gnd WL123 net124 vcc buffer
x225 gnd WL124 net125 vcc buffer
x226 gnd WL125 net126 vcc buffer
x227 gnd WL126 net127 vcc buffer
x228 gnd WL127 net128 vcc buffer
x229 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net129 net130 net131 net132 net133 net134 net135 net136 net137 net138
+ net139 net140 net141 net142 net143 net144 net145 net146 net147 net148 net149 net150 net151 net152 net153
+ net154 net155 net156 net157 net158 net159 net160 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x230 gnd WL128 net129 vcc buffer
x231 gnd WL129 net130 vcc buffer
x232 gnd WL130 net131 vcc buffer
x233 gnd WL131 net132 vcc buffer
x234 gnd WL132 net133 vcc buffer
x235 gnd WL133 net134 vcc buffer
x236 gnd WL134 net135 vcc buffer
x237 gnd WL135 net136 vcc buffer
x238 gnd WL136 net137 vcc buffer
x239 gnd WL137 net138 vcc buffer
x240 gnd WL138 net139 vcc buffer
x241 gnd WL139 net140 vcc buffer
x242 gnd WL140 net141 vcc buffer
x243 gnd WL141 net142 vcc buffer
x244 gnd WL142 net143 vcc buffer
x245 gnd WL143 net144 vcc buffer
x246 gnd WL144 net145 vcc buffer
x247 gnd WL145 net146 vcc buffer
x248 gnd WL146 net147 vcc buffer
x249 gnd WL147 net148 vcc buffer
x250 gnd WL148 net149 vcc buffer
x251 gnd WL149 net150 vcc buffer
x252 gnd WL150 net151 vcc buffer
x253 gnd WL151 net152 vcc buffer
x254 gnd WL152 net153 vcc buffer
x255 gnd WL153 net154 vcc buffer
x256 gnd WL154 net155 vcc buffer
x257 gnd WL155 net156 vcc buffer
x258 gnd WL156 net157 vcc buffer
x259 gnd WL157 net158 vcc buffer
x260 gnd WL158 net159 vcc buffer
x261 gnd WL159 net160 vcc buffer
x262 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net161 net162 net163 net164 net165 net166 net167 net168 net169 net170
+ net171 net172 net173 net174 net175 net176 net177 net178 net179 net180 net181 net182 net183 net184 net185
+ net186 net187 net188 net189 net190 net191 net192 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x263 gnd WL160 net161 vcc buffer
x264 gnd WL161 net162 vcc buffer
x265 gnd WL162 net163 vcc buffer
x266 gnd WL163 net164 vcc buffer
x267 gnd WL164 net165 vcc buffer
x268 gnd WL165 net166 vcc buffer
x269 gnd WL166 net167 vcc buffer
x270 gnd WL167 net168 vcc buffer
x271 gnd WL168 net169 vcc buffer
x272 gnd WL169 net170 vcc buffer
x273 gnd WL170 net171 vcc buffer
x274 gnd WL171 net172 vcc buffer
x275 gnd WL172 net173 vcc buffer
x276 gnd WL173 net174 vcc buffer
x277 gnd WL174 net175 vcc buffer
x278 gnd WL175 net176 vcc buffer
x279 gnd WL176 net177 vcc buffer
x280 gnd WL177 net178 vcc buffer
x281 gnd WL178 net179 vcc buffer
x282 gnd WL179 net180 vcc buffer
x283 gnd WL180 net181 vcc buffer
x284 gnd WL181 net182 vcc buffer
x285 gnd WL182 net183 vcc buffer
x286 gnd WL183 net184 vcc buffer
x287 gnd WL184 net185 vcc buffer
x288 gnd WL185 net186 vcc buffer
x289 gnd WL186 net187 vcc buffer
x290 gnd WL187 net188 vcc buffer
x291 gnd WL188 net189 vcc buffer
x292 gnd WL189 net190 vcc buffer
x293 gnd WL190 net191 vcc buffer
x294 gnd WL191 net192 vcc buffer
x295 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net193 net194 net195 net196 net197 net198 net199 net200 net201 net202
+ net203 net204 net205 net206 net207 net208 net209 net210 net211 net212 net213 net214 net215 net216 net217
+ net218 net219 net220 net221 net222 net223 net224 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x296 gnd WL192 net193 vcc buffer
x297 gnd WL193 net194 vcc buffer
x298 gnd WL194 net195 vcc buffer
x299 gnd WL195 net196 vcc buffer
x300 gnd WL196 net197 vcc buffer
x301 gnd WL197 net198 vcc buffer
x302 gnd WL198 net199 vcc buffer
x303 gnd WL199 net200 vcc buffer
x304 gnd WL200 net201 vcc buffer
x305 gnd WL201 net202 vcc buffer
x306 gnd WL202 net203 vcc buffer
x307 gnd WL203 net204 vcc buffer
x308 gnd WL204 net205 vcc buffer
x309 gnd WL205 net206 vcc buffer
x310 gnd WL206 net207 vcc buffer
x311 gnd WL207 net208 vcc buffer
x312 gnd WL208 net209 vcc buffer
x313 gnd WL209 net210 vcc buffer
x314 gnd WL210 net211 vcc buffer
x315 gnd WL211 net212 vcc buffer
x316 gnd WL212 net213 vcc buffer
x317 gnd WL213 net214 vcc buffer
x318 gnd WL214 net215 vcc buffer
x319 gnd WL215 net216 vcc buffer
x320 gnd WL216 net217 vcc buffer
x321 gnd WL217 net218 vcc buffer
x322 gnd WL218 net219 vcc buffer
x323 gnd WL219 net220 vcc buffer
x324 gnd WL220 net221 vcc buffer
x325 gnd WL221 net222 vcc buffer
x326 gnd WL222 net223 vcc buffer
x327 gnd WL223 net224 vcc buffer
x328 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net225 net226 net227 net228 net229 net230 net231 net232 net233 net234
+ net235 net236 net237 net238 net239 net240 net241 net242 net243 net244 net245 net246 net247 net248 net249
+ net250 net251 net252 net253 net254 net255 net256 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x329 gnd WL224 net225 vcc buffer
x330 gnd WL225 net226 vcc buffer
x331 gnd WL226 net227 vcc buffer
x332 gnd WL227 net228 vcc buffer
x333 gnd WL228 net229 vcc buffer
x334 gnd WL229 net230 vcc buffer
x335 gnd WL230 net231 vcc buffer
x336 gnd WL231 net232 vcc buffer
x337 gnd WL232 net233 vcc buffer
x338 gnd WL233 net234 vcc buffer
x339 gnd WL234 net235 vcc buffer
x340 gnd WL235 net236 vcc buffer
x341 gnd WL236 net237 vcc buffer
x342 gnd WL237 net238 vcc buffer
x343 gnd WL238 net239 vcc buffer
x344 gnd WL239 net240 vcc buffer
x345 gnd WL240 net241 vcc buffer
x346 gnd WL241 net242 vcc buffer
x347 gnd WL242 net243 vcc buffer
x348 gnd WL243 net244 vcc buffer
x349 gnd WL244 net245 vcc buffer
x350 gnd WL245 net246 vcc buffer
x351 gnd WL246 net247 vcc buffer
x352 gnd WL247 net248 vcc buffer
x353 gnd WL248 net249 vcc buffer
x354 gnd WL249 net250 vcc buffer
x355 gnd WL250 net251 vcc buffer
x356 gnd WL251 net252 vcc buffer
x357 gnd WL252 net253 vcc buffer
x358 gnd WL253 net254 vcc buffer
x359 gnd WL254 net255 vcc buffer
x360 gnd WL255 net256 vcc buffer
x361 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net257 net258 net259 net260 net261 net262 net263 net264 net265 net266
+ net267 net268 net269 net270 net271 net272 net273 net274 net275 net276 net277 net278 net279 net280 net281
+ net282 net283 net284 net285 net286 net287 net288 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x362 gnd WL256 net257 vcc buffer
x363 gnd WL257 net258 vcc buffer
x364 gnd WL258 net259 vcc buffer
x365 gnd WL259 net260 vcc buffer
x366 gnd WL260 net261 vcc buffer
x367 gnd WL261 net262 vcc buffer
x368 gnd WL262 net263 vcc buffer
x369 gnd WL263 net264 vcc buffer
x370 gnd WL264 net265 vcc buffer
x371 gnd WL265 net266 vcc buffer
x372 gnd WL266 net267 vcc buffer
x373 gnd WL267 net268 vcc buffer
x374 gnd WL268 net269 vcc buffer
x375 gnd WL269 net270 vcc buffer
x376 gnd WL270 net271 vcc buffer
x377 gnd WL271 net272 vcc buffer
x378 gnd WL272 net273 vcc buffer
x379 gnd WL273 net274 vcc buffer
x380 gnd WL274 net275 vcc buffer
x381 gnd WL275 net276 vcc buffer
x382 gnd WL276 net277 vcc buffer
x383 gnd WL277 net278 vcc buffer
x384 gnd WL278 net279 vcc buffer
x385 gnd WL279 net280 vcc buffer
x386 gnd WL280 net281 vcc buffer
x387 gnd WL281 net282 vcc buffer
x388 gnd WL282 net283 vcc buffer
x389 gnd WL283 net284 vcc buffer
x390 gnd WL284 net285 vcc buffer
x391 gnd WL285 net286 vcc buffer
x392 gnd WL286 net287 vcc buffer
x393 gnd WL287 net288 vcc buffer
x394 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net289 net290 net291 net292 net293 net294 net295 net296 net297 net298
+ net299 net300 net301 net302 net303 net304 net305 net306 net307 net308 net309 net310 net311 net312 net313
+ net314 net315 net316 net317 net318 net319 net320 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x395 gnd WL288 net289 vcc buffer
x396 gnd WL289 net290 vcc buffer
x397 gnd WL290 net291 vcc buffer
x398 gnd WL291 net292 vcc buffer
x399 gnd WL292 net293 vcc buffer
x400 gnd WL293 net294 vcc buffer
x401 gnd WL294 net295 vcc buffer
x402 gnd WL295 net296 vcc buffer
x403 gnd WL296 net297 vcc buffer
x404 gnd WL297 net298 vcc buffer
x405 gnd WL298 net299 vcc buffer
x406 gnd WL299 net300 vcc buffer
x407 gnd WL300 net301 vcc buffer
x408 gnd WL301 net302 vcc buffer
x409 gnd WL302 net303 vcc buffer
x410 gnd WL303 net304 vcc buffer
x411 gnd WL304 net305 vcc buffer
x412 gnd WL305 net306 vcc buffer
x413 gnd WL306 net307 vcc buffer
x414 gnd WL307 net308 vcc buffer
x415 gnd WL308 net309 vcc buffer
x416 gnd WL309 net310 vcc buffer
x417 gnd WL310 net311 vcc buffer
x418 gnd WL311 net312 vcc buffer
x419 gnd WL312 net313 vcc buffer
x420 gnd WL313 net314 vcc buffer
x421 gnd WL314 net315 vcc buffer
x422 gnd WL315 net316 vcc buffer
x423 gnd WL316 net317 vcc buffer
x424 gnd WL317 net318 vcc buffer
x425 gnd WL318 net319 vcc buffer
x426 gnd WL319 net320 vcc buffer
x427 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net321 net322 net323 net324 net325 net326 net327 net328 net329 net330
+ net331 net332 net333 net334 net335 net336 net337 net338 net339 net340 net341 net342 net343 net344 net345
+ net346 net347 net348 net349 net350 net351 net352 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x428 gnd WL320 net321 vcc buffer
x429 gnd WL321 net322 vcc buffer
x430 gnd WL322 net323 vcc buffer
x431 gnd WL323 net324 vcc buffer
x432 gnd WL324 net325 vcc buffer
x433 gnd WL325 net326 vcc buffer
x434 gnd WL326 net327 vcc buffer
x435 gnd WL327 net328 vcc buffer
x436 gnd WL328 net329 vcc buffer
x437 gnd WL329 net330 vcc buffer
x438 gnd WL330 net331 vcc buffer
x439 gnd WL331 net332 vcc buffer
x440 gnd WL332 net333 vcc buffer
x441 gnd WL333 net334 vcc buffer
x442 gnd WL334 net335 vcc buffer
x443 gnd WL335 net336 vcc buffer
x444 gnd WL336 net337 vcc buffer
x445 gnd WL337 net338 vcc buffer
x446 gnd WL338 net339 vcc buffer
x447 gnd WL339 net340 vcc buffer
x448 gnd WL340 net341 vcc buffer
x449 gnd WL341 net342 vcc buffer
x450 gnd WL342 net343 vcc buffer
x451 gnd WL343 net344 vcc buffer
x452 gnd WL344 net345 vcc buffer
x453 gnd WL345 net346 vcc buffer
x454 gnd WL346 net347 vcc buffer
x455 gnd WL347 net348 vcc buffer
x456 gnd WL348 net349 vcc buffer
x457 gnd WL349 net350 vcc buffer
x458 gnd WL350 net351 vcc buffer
x459 gnd WL351 net352 vcc buffer
x460 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net353 net354 net355 net356 net357 net358 net359 net360 net361 net362
+ net363 net364 net365 net366 net367 net368 net369 net370 net371 net372 net373 net374 net375 net376 net377
+ net378 net379 net380 net381 net382 net383 net384 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x461 gnd WL352 net353 vcc buffer
x462 gnd WL353 net354 vcc buffer
x463 gnd WL354 net355 vcc buffer
x464 gnd WL355 net356 vcc buffer
x465 gnd WL356 net357 vcc buffer
x466 gnd WL357 net358 vcc buffer
x467 gnd WL358 net359 vcc buffer
x468 gnd WL359 net360 vcc buffer
x469 gnd WL360 net361 vcc buffer
x470 gnd WL361 net362 vcc buffer
x471 gnd WL362 net363 vcc buffer
x472 gnd WL363 net364 vcc buffer
x473 gnd WL364 net365 vcc buffer
x474 gnd WL365 net366 vcc buffer
x475 gnd WL366 net367 vcc buffer
x476 gnd WL367 net368 vcc buffer
x477 gnd WL368 net369 vcc buffer
x478 gnd WL369 net370 vcc buffer
x479 gnd WL370 net371 vcc buffer
x480 gnd WL371 net372 vcc buffer
x481 gnd WL372 net373 vcc buffer
x482 gnd WL373 net374 vcc buffer
x483 gnd WL374 net375 vcc buffer
x484 gnd WL375 net376 vcc buffer
x485 gnd WL376 net377 vcc buffer
x486 gnd WL377 net378 vcc buffer
x487 gnd WL378 net379 vcc buffer
x488 gnd WL379 net380 vcc buffer
x489 gnd WL380 net381 vcc buffer
x490 gnd WL381 net382 vcc buffer
x491 gnd WL382 net383 vcc buffer
x492 gnd WL383 net384 vcc buffer
x493 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net385 net386 net387 net388 net389 net390 net391 net392 net393 net394
+ net395 net396 net397 net398 net399 net400 net401 net402 net403 net404 net405 net406 net407 net408 net409
+ net410 net411 net412 net413 net414 net415 net416 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x494 gnd WL384 net385 vcc buffer
x495 gnd WL385 net386 vcc buffer
x496 gnd WL386 net387 vcc buffer
x497 gnd WL387 net388 vcc buffer
x498 gnd WL388 net389 vcc buffer
x499 gnd WL389 net390 vcc buffer
x500 gnd WL390 net391 vcc buffer
x501 gnd WL391 net392 vcc buffer
x502 gnd WL392 net393 vcc buffer
x503 gnd WL393 net394 vcc buffer
x504 gnd WL394 net395 vcc buffer
x505 gnd WL395 net396 vcc buffer
x506 gnd WL396 net397 vcc buffer
x507 gnd WL397 net398 vcc buffer
x508 gnd WL398 net399 vcc buffer
x509 gnd WL399 net400 vcc buffer
x510 gnd WL400 net401 vcc buffer
x511 gnd WL401 net402 vcc buffer
x512 gnd WL402 net403 vcc buffer
x513 gnd WL403 net404 vcc buffer
x514 gnd WL404 net405 vcc buffer
x515 gnd WL405 net406 vcc buffer
x516 gnd WL406 net407 vcc buffer
x517 gnd WL407 net408 vcc buffer
x518 gnd WL408 net409 vcc buffer
x519 gnd WL409 net410 vcc buffer
x520 gnd WL410 net411 vcc buffer
x521 gnd WL411 net412 vcc buffer
x522 gnd WL412 net413 vcc buffer
x523 gnd WL413 net414 vcc buffer
x524 gnd WL414 net415 vcc buffer
x525 gnd WL415 net416 vcc buffer
x526 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net417 net418 net419 net420 net421 net422 net423 net424 net425 net426
+ net427 net428 net429 net430 net431 net432 net433 net434 net435 net436 net437 net438 net439 net440 net441
+ net442 net443 net444 net445 net446 net447 net448 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x527 gnd WL416 net417 vcc buffer
x528 gnd WL417 net418 vcc buffer
x529 gnd WL418 net419 vcc buffer
x530 gnd WL419 net420 vcc buffer
x531 gnd WL420 net421 vcc buffer
x532 gnd WL421 net422 vcc buffer
x533 gnd WL422 net423 vcc buffer
x534 gnd WL423 net424 vcc buffer
x535 gnd WL424 net425 vcc buffer
x536 gnd WL425 net426 vcc buffer
x537 gnd WL426 net427 vcc buffer
x538 gnd WL427 net428 vcc buffer
x539 gnd WL428 net429 vcc buffer
x540 gnd WL429 net430 vcc buffer
x541 gnd WL430 net431 vcc buffer
x542 gnd WL431 net432 vcc buffer
x543 gnd WL432 net433 vcc buffer
x544 gnd WL433 net434 vcc buffer
x545 gnd WL434 net435 vcc buffer
x546 gnd WL435 net436 vcc buffer
x547 gnd WL436 net437 vcc buffer
x548 gnd WL437 net438 vcc buffer
x549 gnd WL438 net439 vcc buffer
x550 gnd WL439 net440 vcc buffer
x551 gnd WL440 net441 vcc buffer
x552 gnd WL441 net442 vcc buffer
x553 gnd WL442 net443 vcc buffer
x554 gnd WL443 net444 vcc buffer
x555 gnd WL444 net445 vcc buffer
x556 gnd WL445 net446 vcc buffer
x557 gnd WL446 net447 vcc buffer
x558 gnd WL447 net448 vcc buffer
x559 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net449 net450 net451 net452 net453 net454 net455 net456 net457 net458
+ net459 net460 net461 net462 net463 net464 net465 net466 net467 net468 net469 net470 net471 net472 net473
+ net474 net475 net476 net477 net478 net479 net480 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x560 gnd WL448 net449 vcc buffer
x561 gnd WL449 net450 vcc buffer
x562 gnd WL450 net451 vcc buffer
x563 gnd WL451 net452 vcc buffer
x564 gnd WL452 net453 vcc buffer
x565 gnd WL453 net454 vcc buffer
x566 gnd WL454 net455 vcc buffer
x567 gnd WL455 net456 vcc buffer
x568 gnd WL456 net457 vcc buffer
x569 gnd WL457 net458 vcc buffer
x570 gnd WL458 net459 vcc buffer
x571 gnd WL459 net460 vcc buffer
x572 gnd WL460 net461 vcc buffer
x573 gnd WL461 net462 vcc buffer
x574 gnd WL462 net463 vcc buffer
x575 gnd WL463 net464 vcc buffer
x576 gnd WL464 net465 vcc buffer
x577 gnd WL465 net466 vcc buffer
x578 gnd WL466 net467 vcc buffer
x579 gnd WL467 net468 vcc buffer
x580 gnd WL468 net469 vcc buffer
x581 gnd WL469 net470 vcc buffer
x582 gnd WL470 net471 vcc buffer
x583 gnd WL471 net472 vcc buffer
x584 gnd WL472 net473 vcc buffer
x585 gnd WL473 net474 vcc buffer
x586 gnd WL474 net475 vcc buffer
x587 gnd WL475 net476 vcc buffer
x588 gnd WL476 net477 vcc buffer
x589 gnd WL477 net478 vcc buffer
x590 gnd WL478 net479 vcc buffer
x591 gnd WL479 net480 vcc buffer
x592 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net481 net482 net483 net484 net485 net486 net487 net488 net489 net490
+ net491 net492 net493 net494 net495 net496 net497 net498 net499 net500 net501 net502 net503 net504 net505
+ net506 net507 net508 net509 net510 net511 net512 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x593 gnd WL480 net481 vcc buffer
x594 gnd WL481 net482 vcc buffer
x595 gnd WL482 net483 vcc buffer
x596 gnd WL483 net484 vcc buffer
x597 gnd WL484 net485 vcc buffer
x598 gnd WL485 net486 vcc buffer
x599 gnd WL486 net487 vcc buffer
x600 gnd WL487 net488 vcc buffer
x601 gnd WL488 net489 vcc buffer
x602 gnd WL489 net490 vcc buffer
x603 gnd WL490 net491 vcc buffer
x604 gnd WL491 net492 vcc buffer
x605 gnd WL492 net493 vcc buffer
x606 gnd WL493 net494 vcc buffer
x607 gnd WL494 net495 vcc buffer
x608 gnd WL495 net496 vcc buffer
x609 gnd WL496 net497 vcc buffer
x610 gnd WL497 net498 vcc buffer
x611 gnd WL498 net499 vcc buffer
x612 gnd WL499 net500 vcc buffer
x613 gnd WL500 net501 vcc buffer
x614 gnd WL501 net502 vcc buffer
x615 gnd WL502 net503 vcc buffer
x616 gnd WL503 net504 vcc buffer
x617 gnd WL504 net505 vcc buffer
x618 gnd WL505 net506 vcc buffer
x619 gnd WL506 net507 vcc buffer
x620 gnd WL507 net508 vcc buffer
x621 gnd WL508 net509 vcc buffer
x622 gnd WL509 net510 vcc buffer
x623 gnd WL510 net511 vcc buffer
x624 gnd WL511 net512 vcc buffer
x625 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net513 net514 net515 net516 net517 net518 net519 net520 net521 net522
+ net523 net524 net525 net526 net527 net528 net529 net530 net531 net532 net533 net534 net535 net536 net537
+ net538 net539 net540 net541 net542 net543 net544 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x626 gnd WL512 net513 vcc buffer
x627 gnd WL513 net514 vcc buffer
x628 gnd WL514 net515 vcc buffer
x629 gnd WL515 net516 vcc buffer
x630 gnd WL516 net517 vcc buffer
x631 gnd WL517 net518 vcc buffer
x632 gnd WL518 net519 vcc buffer
x633 gnd WL519 net520 vcc buffer
x634 gnd WL520 net521 vcc buffer
x635 gnd WL521 net522 vcc buffer
x636 gnd WL522 net523 vcc buffer
x637 gnd WL523 net524 vcc buffer
x638 gnd WL524 net525 vcc buffer
x639 gnd WL525 net526 vcc buffer
x640 gnd WL526 net527 vcc buffer
x641 gnd WL527 net528 vcc buffer
x642 gnd WL528 net529 vcc buffer
x643 gnd WL529 net530 vcc buffer
x644 gnd WL530 net531 vcc buffer
x645 gnd WL531 net532 vcc buffer
x646 gnd WL532 net533 vcc buffer
x647 gnd WL533 net534 vcc buffer
x648 gnd WL534 net535 vcc buffer
x649 gnd WL535 net536 vcc buffer
x650 gnd WL536 net537 vcc buffer
x651 gnd WL537 net538 vcc buffer
x652 gnd WL538 net539 vcc buffer
x653 gnd WL539 net540 vcc buffer
x654 gnd WL540 net541 vcc buffer
x655 gnd WL541 net542 vcc buffer
x656 gnd WL542 net543 vcc buffer
x657 gnd WL543 net544 vcc buffer
x658 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net545 net546 net547 net548 net549 net550 net551 net552 net553 net554
+ net555 net556 net557 net558 net559 net560 net561 net562 net563 net564 net565 net566 net567 net568 net569
+ net570 net571 net572 net573 net574 net575 net576 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x659 gnd WL544 net545 vcc buffer
x660 gnd WL545 net546 vcc buffer
x661 gnd WL546 net547 vcc buffer
x662 gnd WL547 net548 vcc buffer
x663 gnd WL548 net549 vcc buffer
x664 gnd WL549 net550 vcc buffer
x665 gnd WL550 net551 vcc buffer
x666 gnd WL551 net552 vcc buffer
x667 gnd WL552 net553 vcc buffer
x668 gnd WL553 net554 vcc buffer
x669 gnd WL554 net555 vcc buffer
x670 gnd WL555 net556 vcc buffer
x671 gnd WL556 net557 vcc buffer
x672 gnd WL557 net558 vcc buffer
x673 gnd WL558 net559 vcc buffer
x674 gnd WL559 net560 vcc buffer
x675 gnd WL560 net561 vcc buffer
x676 gnd WL561 net562 vcc buffer
x677 gnd WL562 net563 vcc buffer
x678 gnd WL563 net564 vcc buffer
x679 gnd WL564 net565 vcc buffer
x680 gnd WL565 net566 vcc buffer
x681 gnd WL566 net567 vcc buffer
x682 gnd WL567 net568 vcc buffer
x683 gnd WL568 net569 vcc buffer
x684 gnd WL569 net570 vcc buffer
x685 gnd WL570 net571 vcc buffer
x686 gnd WL571 net572 vcc buffer
x687 gnd WL572 net573 vcc buffer
x688 gnd WL573 net574 vcc buffer
x689 gnd WL574 net575 vcc buffer
x690 gnd WL575 net576 vcc buffer
x691 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net577 net578 net579 net580 net581 net582 net583 net584 net585 net586
+ net587 net588 net589 net590 net591 net592 net593 net594 net595 net596 net597 net598 net599 net600 net601
+ net602 net603 net604 net605 net606 net607 net608 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x692 gnd WL576 net577 vcc buffer
x693 gnd WL577 net578 vcc buffer
x694 gnd WL578 net579 vcc buffer
x695 gnd WL579 net580 vcc buffer
x696 gnd WL580 net581 vcc buffer
x697 gnd WL581 net582 vcc buffer
x698 gnd WL582 net583 vcc buffer
x699 gnd WL583 net584 vcc buffer
x700 gnd WL584 net585 vcc buffer
x701 gnd WL585 net586 vcc buffer
x702 gnd WL586 net587 vcc buffer
x703 gnd WL587 net588 vcc buffer
x704 gnd WL588 net589 vcc buffer
x705 gnd WL589 net590 vcc buffer
x706 gnd WL590 net591 vcc buffer
x707 gnd WL591 net592 vcc buffer
x708 gnd WL592 net593 vcc buffer
x709 gnd WL593 net594 vcc buffer
x710 gnd WL594 net595 vcc buffer
x711 gnd WL595 net596 vcc buffer
x712 gnd WL596 net597 vcc buffer
x713 gnd WL597 net598 vcc buffer
x714 gnd WL598 net599 vcc buffer
x715 gnd WL599 net600 vcc buffer
x716 gnd WL600 net601 vcc buffer
x717 gnd WL601 net602 vcc buffer
x718 gnd WL602 net603 vcc buffer
x719 gnd WL603 net604 vcc buffer
x720 gnd WL604 net605 vcc buffer
x721 gnd WL605 net606 vcc buffer
x722 gnd WL606 net607 vcc buffer
x723 gnd WL607 net608 vcc buffer
x724 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net609 net610 net611 net612 net613 net614 net615 net616 net617 net618
+ net619 net620 net621 net622 net623 net624 net625 net626 net627 net628 net629 net630 net631 net632 net633
+ net634 net635 net636 net637 net638 net639 net640 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x725 gnd WL608 net609 vcc buffer
x726 gnd WL609 net610 vcc buffer
x727 gnd WL610 net611 vcc buffer
x728 gnd WL611 net612 vcc buffer
x729 gnd WL612 net613 vcc buffer
x730 gnd WL613 net614 vcc buffer
x731 gnd WL614 net615 vcc buffer
x732 gnd WL615 net616 vcc buffer
x733 gnd WL616 net617 vcc buffer
x734 gnd WL617 net618 vcc buffer
x735 gnd WL618 net619 vcc buffer
x736 gnd WL619 net620 vcc buffer
x737 gnd WL620 net621 vcc buffer
x738 gnd WL621 net622 vcc buffer
x739 gnd WL622 net623 vcc buffer
x740 gnd WL623 net624 vcc buffer
x741 gnd WL624 net625 vcc buffer
x742 gnd WL625 net626 vcc buffer
x743 gnd WL626 net627 vcc buffer
x744 gnd WL627 net628 vcc buffer
x745 gnd WL628 net629 vcc buffer
x746 gnd WL629 net630 vcc buffer
x747 gnd WL630 net631 vcc buffer
x748 gnd WL631 net632 vcc buffer
x749 gnd WL632 net633 vcc buffer
x750 gnd WL633 net634 vcc buffer
x751 gnd WL634 net635 vcc buffer
x752 gnd WL635 net636 vcc buffer
x753 gnd WL636 net637 vcc buffer
x754 gnd WL637 net638 vcc buffer
x755 gnd WL638 net639 vcc buffer
x756 gnd WL639 net640 vcc buffer
x757 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net641 net642 net643 net644 net645 net646 net647 net648 net649 net650
+ net651 net652 net653 net654 net655 net656 net657 net658 net659 net660 net661 net662 net663 net664 net665
+ net666 net667 net668 net669 net670 net671 net672 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x758 gnd WL640 net641 vcc buffer
x759 gnd WL641 net642 vcc buffer
x760 gnd WL642 net643 vcc buffer
x761 gnd WL643 net644 vcc buffer
x762 gnd WL644 net645 vcc buffer
x763 gnd WL645 net646 vcc buffer
x764 gnd WL646 net647 vcc buffer
x765 gnd WL647 net648 vcc buffer
x766 gnd WL648 net649 vcc buffer
x767 gnd WL649 net650 vcc buffer
x768 gnd WL650 net651 vcc buffer
x769 gnd WL651 net652 vcc buffer
x770 gnd WL652 net653 vcc buffer
x771 gnd WL653 net654 vcc buffer
x772 gnd WL654 net655 vcc buffer
x773 gnd WL655 net656 vcc buffer
x774 gnd WL656 net657 vcc buffer
x775 gnd WL657 net658 vcc buffer
x776 gnd WL658 net659 vcc buffer
x777 gnd WL659 net660 vcc buffer
x778 gnd WL660 net661 vcc buffer
x779 gnd WL661 net662 vcc buffer
x780 gnd WL662 net663 vcc buffer
x781 gnd WL663 net664 vcc buffer
x782 gnd WL664 net665 vcc buffer
x783 gnd WL665 net666 vcc buffer
x784 gnd WL666 net667 vcc buffer
x785 gnd WL667 net668 vcc buffer
x786 gnd WL668 net669 vcc buffer
x787 gnd WL669 net670 vcc buffer
x788 gnd WL670 net671 vcc buffer
x789 gnd WL671 net672 vcc buffer
x790 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net673 net674 net675 net676 net677 net678 net679 net680 net681 net682
+ net683 net684 net685 net686 net687 net688 net689 net690 net691 net692 net693 net694 net695 net696 net697
+ net698 net699 net700 net701 net702 net703 net704 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x791 gnd WL672 net673 vcc buffer
x792 gnd WL673 net674 vcc buffer
x793 gnd WL674 net675 vcc buffer
x794 gnd WL675 net676 vcc buffer
x795 gnd WL676 net677 vcc buffer
x796 gnd WL677 net678 vcc buffer
x797 gnd WL678 net679 vcc buffer
x798 gnd WL679 net680 vcc buffer
x799 gnd WL680 net681 vcc buffer
x800 gnd WL681 net682 vcc buffer
x801 gnd WL682 net683 vcc buffer
x802 gnd WL683 net684 vcc buffer
x803 gnd WL684 net685 vcc buffer
x804 gnd WL685 net686 vcc buffer
x805 gnd WL686 net687 vcc buffer
x806 gnd WL687 net688 vcc buffer
x807 gnd WL688 net689 vcc buffer
x808 gnd WL689 net690 vcc buffer
x809 gnd WL690 net691 vcc buffer
x810 gnd WL691 net692 vcc buffer
x811 gnd WL692 net693 vcc buffer
x812 gnd WL693 net694 vcc buffer
x813 gnd WL694 net695 vcc buffer
x814 gnd WL695 net696 vcc buffer
x815 gnd WL696 net697 vcc buffer
x816 gnd WL697 net698 vcc buffer
x817 gnd WL698 net699 vcc buffer
x818 gnd WL699 net700 vcc buffer
x819 gnd WL700 net701 vcc buffer
x820 gnd WL701 net702 vcc buffer
x821 gnd WL702 net703 vcc buffer
x822 gnd WL703 net704 vcc buffer
x823 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net705 net706 net707 net708 net709 net710 net711 net712 net713 net714
+ net715 net716 net717 net718 net719 net720 net721 net722 net723 net724 net725 net726 net727 net728 net729
+ net730 net731 net732 net733 net734 net735 net736 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x824 gnd WL704 net705 vcc buffer
x825 gnd WL705 net706 vcc buffer
x826 gnd WL706 net707 vcc buffer
x827 gnd WL707 net708 vcc buffer
x828 gnd WL708 net709 vcc buffer
x829 gnd WL709 net710 vcc buffer
x830 gnd WL710 net711 vcc buffer
x831 gnd WL711 net712 vcc buffer
x832 gnd WL712 net713 vcc buffer
x833 gnd WL713 net714 vcc buffer
x834 gnd WL714 net715 vcc buffer
x835 gnd WL715 net716 vcc buffer
x836 gnd WL716 net717 vcc buffer
x837 gnd WL717 net718 vcc buffer
x838 gnd WL718 net719 vcc buffer
x839 gnd WL719 net720 vcc buffer
x840 gnd WL720 net721 vcc buffer
x841 gnd WL721 net722 vcc buffer
x842 gnd WL722 net723 vcc buffer
x843 gnd WL723 net724 vcc buffer
x844 gnd WL724 net725 vcc buffer
x845 gnd WL725 net726 vcc buffer
x846 gnd WL726 net727 vcc buffer
x847 gnd WL727 net728 vcc buffer
x848 gnd WL728 net729 vcc buffer
x849 gnd WL729 net730 vcc buffer
x850 gnd WL730 net731 vcc buffer
x851 gnd WL731 net732 vcc buffer
x852 gnd WL732 net733 vcc buffer
x853 gnd WL733 net734 vcc buffer
x854 gnd WL734 net735 vcc buffer
x855 gnd WL735 net736 vcc buffer
x856 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net737 net738 net739 net740 net741 net742 net743 net744 net745 net746
+ net747 net748 net749 net750 net751 net752 net753 net754 net755 net756 net757 net758 net759 net760 net761
+ net762 net763 net764 net765 net766 net767 net768 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x857 gnd WL736 net737 vcc buffer
x858 gnd WL737 net738 vcc buffer
x859 gnd WL738 net739 vcc buffer
x860 gnd WL739 net740 vcc buffer
x861 gnd WL740 net741 vcc buffer
x862 gnd WL741 net742 vcc buffer
x863 gnd WL742 net743 vcc buffer
x864 gnd WL743 net744 vcc buffer
x865 gnd WL744 net745 vcc buffer
x866 gnd WL745 net746 vcc buffer
x867 gnd WL746 net747 vcc buffer
x868 gnd WL747 net748 vcc buffer
x869 gnd WL748 net749 vcc buffer
x870 gnd WL749 net750 vcc buffer
x871 gnd WL750 net751 vcc buffer
x872 gnd WL751 net752 vcc buffer
x873 gnd WL752 net753 vcc buffer
x874 gnd WL753 net754 vcc buffer
x875 gnd WL754 net755 vcc buffer
x876 gnd WL755 net756 vcc buffer
x877 gnd WL756 net757 vcc buffer
x878 gnd WL757 net758 vcc buffer
x879 gnd WL758 net759 vcc buffer
x880 gnd WL759 net760 vcc buffer
x881 gnd WL760 net761 vcc buffer
x882 gnd WL761 net762 vcc buffer
x883 gnd WL762 net763 vcc buffer
x884 gnd WL763 net764 vcc buffer
x885 gnd WL764 net765 vcc buffer
x886 gnd WL765 net766 vcc buffer
x887 gnd WL766 net767 vcc buffer
x888 gnd WL767 net768 vcc buffer
x889 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net769 net770 net771 net772 net773 net774 net775 net776 net777 net778
+ net779 net780 net781 net782 net783 net784 net785 net786 net787 net788 net789 net790 net791 net792 net793
+ net794 net795 net796 net797 net798 net799 net800 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x890 gnd WL768 net769 vcc buffer
x891 gnd WL769 net770 vcc buffer
x892 gnd WL770 net771 vcc buffer
x893 gnd WL771 net772 vcc buffer
x894 gnd WL772 net773 vcc buffer
x895 gnd WL773 net774 vcc buffer
x896 gnd WL774 net775 vcc buffer
x897 gnd WL775 net776 vcc buffer
x898 gnd WL776 net777 vcc buffer
x899 gnd WL777 net778 vcc buffer
x900 gnd WL778 net779 vcc buffer
x901 gnd WL779 net780 vcc buffer
x902 gnd WL780 net781 vcc buffer
x903 gnd WL781 net782 vcc buffer
x904 gnd WL782 net783 vcc buffer
x905 gnd WL783 net784 vcc buffer
x906 gnd WL784 net785 vcc buffer
x907 gnd WL785 net786 vcc buffer
x908 gnd WL786 net787 vcc buffer
x909 gnd WL787 net788 vcc buffer
x910 gnd WL788 net789 vcc buffer
x911 gnd WL789 net790 vcc buffer
x912 gnd WL790 net791 vcc buffer
x913 gnd WL791 net792 vcc buffer
x914 gnd WL792 net793 vcc buffer
x915 gnd WL793 net794 vcc buffer
x916 gnd WL794 net795 vcc buffer
x917 gnd WL795 net796 vcc buffer
x918 gnd WL796 net797 vcc buffer
x919 gnd WL797 net798 vcc buffer
x920 gnd WL798 net799 vcc buffer
x921 gnd WL799 net800 vcc buffer
x922 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net801 net802 net803 net804 net805 net806 net807 net808 net809 net810
+ net811 net812 net813 net814 net815 net816 net817 net818 net819 net820 net821 net822 net823 net824 net825
+ net826 net827 net828 net829 net830 net831 net832 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x923 gnd WL800 net801 vcc buffer
x924 gnd WL801 net802 vcc buffer
x925 gnd WL802 net803 vcc buffer
x926 gnd WL803 net804 vcc buffer
x927 gnd WL804 net805 vcc buffer
x928 gnd WL805 net806 vcc buffer
x929 gnd WL806 net807 vcc buffer
x930 gnd WL807 net808 vcc buffer
x931 gnd WL808 net809 vcc buffer
x932 gnd WL809 net810 vcc buffer
x933 gnd WL810 net811 vcc buffer
x934 gnd WL811 net812 vcc buffer
x935 gnd WL812 net813 vcc buffer
x936 gnd WL813 net814 vcc buffer
x937 gnd WL814 net815 vcc buffer
x938 gnd WL815 net816 vcc buffer
x939 gnd WL816 net817 vcc buffer
x940 gnd WL817 net818 vcc buffer
x941 gnd WL818 net819 vcc buffer
x942 gnd WL819 net820 vcc buffer
x943 gnd WL820 net821 vcc buffer
x944 gnd WL821 net822 vcc buffer
x945 gnd WL822 net823 vcc buffer
x946 gnd WL823 net824 vcc buffer
x947 gnd WL824 net825 vcc buffer
x948 gnd WL825 net826 vcc buffer
x949 gnd WL826 net827 vcc buffer
x950 gnd WL827 net828 vcc buffer
x951 gnd WL828 net829 vcc buffer
x952 gnd WL829 net830 vcc buffer
x953 gnd WL830 net831 vcc buffer
x954 gnd WL831 net832 vcc buffer
x955 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net833 net834 net835 net836 net837 net838 net839 net840 net841 net842
+ net843 net844 net845 net846 net847 net848 net849 net850 net851 net852 net853 net854 net855 net856 net857
+ net858 net859 net860 net861 net862 net863 net864 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x956 gnd WL832 net833 vcc buffer
x957 gnd WL833 net834 vcc buffer
x958 gnd WL834 net835 vcc buffer
x959 gnd WL835 net836 vcc buffer
x960 gnd WL836 net837 vcc buffer
x961 gnd WL837 net838 vcc buffer
x962 gnd WL838 net839 vcc buffer
x963 gnd WL839 net840 vcc buffer
x964 gnd WL840 net841 vcc buffer
x965 gnd WL841 net842 vcc buffer
x966 gnd WL842 net843 vcc buffer
x967 gnd WL843 net844 vcc buffer
x968 gnd WL844 net845 vcc buffer
x969 gnd WL845 net846 vcc buffer
x970 gnd WL846 net847 vcc buffer
x971 gnd WL847 net848 vcc buffer
x972 gnd WL848 net849 vcc buffer
x973 gnd WL849 net850 vcc buffer
x974 gnd WL850 net851 vcc buffer
x975 gnd WL851 net852 vcc buffer
x976 gnd WL852 net853 vcc buffer
x977 gnd WL853 net854 vcc buffer
x978 gnd WL854 net855 vcc buffer
x979 gnd WL855 net856 vcc buffer
x980 gnd WL856 net857 vcc buffer
x981 gnd WL857 net858 vcc buffer
x982 gnd WL858 net859 vcc buffer
x983 gnd WL859 net860 vcc buffer
x984 gnd WL860 net861 vcc buffer
x985 gnd WL861 net862 vcc buffer
x986 gnd WL862 net863 vcc buffer
x987 gnd WL863 net864 vcc buffer
x988 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net865 net866 net867 net868 net869 net870 net871 net872 net873 net874
+ net875 net876 net877 net878 net879 net880 net881 net882 net883 net884 net885 net886 net887 net888 net889
+ net890 net891 net892 net893 net894 net895 net896 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x989 gnd WL864 net865 vcc buffer
x990 gnd WL865 net866 vcc buffer
x991 gnd WL866 net867 vcc buffer
x992 gnd WL867 net868 vcc buffer
x993 gnd WL868 net869 vcc buffer
x994 gnd WL869 net870 vcc buffer
x995 gnd WL870 net871 vcc buffer
x996 gnd WL871 net872 vcc buffer
x997 gnd WL872 net873 vcc buffer
x998 gnd WL873 net874 vcc buffer
x999 gnd WL874 net875 vcc buffer
x1000 gnd WL875 net876 vcc buffer
x1001 gnd WL876 net877 vcc buffer
x1002 gnd WL877 net878 vcc buffer
x1003 gnd WL878 net879 vcc buffer
x1004 gnd WL879 net880 vcc buffer
x1005 gnd WL880 net881 vcc buffer
x1006 gnd WL881 net882 vcc buffer
x1007 gnd WL882 net883 vcc buffer
x1008 gnd WL883 net884 vcc buffer
x1009 gnd WL884 net885 vcc buffer
x1010 gnd WL885 net886 vcc buffer
x1011 gnd WL886 net887 vcc buffer
x1012 gnd WL887 net888 vcc buffer
x1013 gnd WL888 net889 vcc buffer
x1014 gnd WL889 net890 vcc buffer
x1015 gnd WL890 net891 vcc buffer
x1016 gnd WL891 net892 vcc buffer
x1017 gnd WL892 net893 vcc buffer
x1018 gnd WL893 net894 vcc buffer
x1019 gnd WL894 net895 vcc buffer
x1020 gnd WL895 net896 vcc buffer
x1021 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5
+ gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net897 net898 net899 net900 net901 net902 net903 net904 net905 net906
+ net907 net908 net909 net910 net911 net912 net913 net914 net915 net916 net917 net918 net919 net920 net921
+ net922 net923 net924 net925 net926 net927 net928 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x1022 gnd WL896 net897 vcc buffer
x1023 gnd WL897 net898 vcc buffer
x1024 gnd WL898 net899 vcc buffer
x1025 gnd WL899 net900 vcc buffer
x1026 gnd WL900 net901 vcc buffer
x1027 gnd WL901 net902 vcc buffer
x1028 gnd WL902 net903 vcc buffer
x1029 gnd WL903 net904 vcc buffer
x1030 gnd WL904 net905 vcc buffer
x1031 gnd WL905 net906 vcc buffer
x1032 gnd WL906 net907 vcc buffer
x1033 gnd WL907 net908 vcc buffer
x1034 gnd WL908 net909 vcc buffer
x1035 gnd WL909 net910 vcc buffer
x1036 gnd WL910 net911 vcc buffer
x1037 gnd WL911 net912 vcc buffer
x1038 gnd WL912 net913 vcc buffer
x1039 gnd WL913 net914 vcc buffer
x1040 gnd WL914 net915 vcc buffer
x1041 gnd WL915 net916 vcc buffer
x1042 gnd WL916 net917 vcc buffer
x1043 gnd WL917 net918 vcc buffer
x1044 gnd WL918 net919 vcc buffer
x1045 gnd WL919 net920 vcc buffer
x1046 gnd WL920 net921 vcc buffer
x1047 gnd WL921 net922 vcc buffer
x1048 gnd WL922 net923 vcc buffer
x1049 gnd WL923 net924 vcc buffer
x1050 gnd WL924 net925 vcc buffer
x1051 gnd WL925 net926 vcc buffer
x1052 gnd WL926 net927 vcc buffer
x1053 gnd WL927 net928 vcc buffer
x1054 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5
+ gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net929 net930 net931 net932 net933 net934 net935 net936 net937 net938
+ net939 net940 net941 net942 net943 net944 net945 net946 net947 net948 net949 net950 net951 net952 net953
+ net954 net955 net956 net957 net958 net959 net960 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x1055 gnd WL928 net929 vcc buffer
x1056 gnd WL929 net930 vcc buffer
x1057 gnd WL930 net931 vcc buffer
x1058 gnd WL931 net932 vcc buffer
x1059 gnd WL932 net933 vcc buffer
x1060 gnd WL933 net934 vcc buffer
x1061 gnd WL934 net935 vcc buffer
x1062 gnd WL935 net936 vcc buffer
x1063 gnd WL936 net937 vcc buffer
x1064 gnd WL937 net938 vcc buffer
x1065 gnd WL938 net939 vcc buffer
x1066 gnd WL939 net940 vcc buffer
x1067 gnd WL940 net941 vcc buffer
x1068 gnd WL941 net942 vcc buffer
x1069 gnd WL942 net943 vcc buffer
x1070 gnd WL943 net944 vcc buffer
x1071 gnd WL944 net945 vcc buffer
x1072 gnd WL945 net946 vcc buffer
x1073 gnd WL946 net947 vcc buffer
x1074 gnd WL947 net948 vcc buffer
x1075 gnd WL948 net949 vcc buffer
x1076 gnd WL949 net950 vcc buffer
x1077 gnd WL950 net951 vcc buffer
x1078 gnd WL951 net952 vcc buffer
x1079 gnd WL952 net953 vcc buffer
x1080 gnd WL953 net954 vcc buffer
x1081 gnd WL954 net955 vcc buffer
x1082 gnd WL955 net956 vcc buffer
x1083 gnd WL956 net957 vcc buffer
x1084 gnd WL957 net958 vcc buffer
x1085 gnd WL958 net959 vcc buffer
x1086 gnd WL959 net960 vcc buffer
x1087 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5
+ gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net961 net962 net963 net964 net965 net966 net967 net968 net969 net970
+ net971 net972 net973 net974 net975 net976 net977 net978 net979 net980 net981 net982 net983 net984 net985
+ net986 net987 net988 net989 net990 net991 net992 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31
+ Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23
+ Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25
+ Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd 32x32_truncation_sram
x1088 gnd WL960 net961 vcc buffer
x1089 gnd WL961 net962 vcc buffer
x1090 gnd WL962 net963 vcc buffer
x1091 gnd WL963 net964 vcc buffer
x1092 gnd WL964 net965 vcc buffer
x1093 gnd WL965 net966 vcc buffer
x1094 gnd WL966 net967 vcc buffer
x1095 gnd WL967 net968 vcc buffer
x1096 gnd WL968 net969 vcc buffer
x1097 gnd WL969 net970 vcc buffer
x1098 gnd WL970 net971 vcc buffer
x1099 gnd WL971 net972 vcc buffer
x1100 gnd WL972 net973 vcc buffer
x1101 gnd WL973 net974 vcc buffer
x1102 gnd WL974 net975 vcc buffer
x1103 gnd WL975 net976 vcc buffer
x1104 gnd WL976 net977 vcc buffer
x1105 gnd WL977 net978 vcc buffer
x1106 gnd WL978 net979 vcc buffer
x1107 gnd WL979 net980 vcc buffer
x1108 gnd WL980 net981 vcc buffer
x1109 gnd WL981 net982 vcc buffer
x1110 gnd WL982 net983 vcc buffer
x1111 gnd WL983 net984 vcc buffer
x1112 gnd WL984 net985 vcc buffer
x1113 gnd WL985 net986 vcc buffer
x1114 gnd WL986 net987 vcc buffer
x1115 gnd WL987 net988 vcc buffer
x1116 gnd WL988 net989 vcc buffer
x1117 gnd WL989 net990 vcc buffer
x1118 gnd WL990 net991 vcc buffer
x1119 gnd WL991 net992 vcc buffer
x1120 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5
+ gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17
+ vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23
+ vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29
+ vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 net993 net994 net995 net996 net997 net998 net999 net1000 net1001 net1002
+ net1003 net1004 net1005 net1006 net1007 net1008 net1009 net1010 net1011 net1012 net1013 net1014 net1015
+ net1016 net1017 net1018 net1019 net1020 net1021 net1022 net1023 net1024 Blb13 Bl13 Blb12 Blb11 Bl11 Blb10
+ Blb9 Bl9 Blb8 Bl8 Blb31 Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10 Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24
+ Bl14 Blb3 Blb23 Bl23 Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19 Blb18 B21 Blb1 Bl22 Bl18 Blb17 Bl17
+ Bl24 Blb16 Bl25 Blb25 Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30 Blb14 Bl1 Blb0 Bl0 gnd
+ 32x32_truncation_sram
x1121 gnd WL992 net993 vcc buffer
x1122 gnd WL993 net994 vcc buffer
x1123 gnd WL994 net995 vcc buffer
x1124 gnd WL995 net996 vcc buffer
x1125 gnd WL996 net997 vcc buffer
x1126 gnd WL997 net998 vcc buffer
x1127 gnd WL998 net999 vcc buffer
x1128 gnd WL999 net1000 vcc buffer
x1129 gnd WL1000 net1001 vcc buffer
x1130 gnd WL1001 net1002 vcc buffer
x1131 gnd WL1002 net1003 vcc buffer
x1132 gnd WL1003 net1004 vcc buffer
x1133 gnd WL1004 net1005 vcc buffer
x1134 gnd WL1005 net1006 vcc buffer
x1135 gnd WL1006 net1007 vcc buffer
x1136 gnd WL1007 net1008 vcc buffer
x1137 gnd WL1008 net1009 vcc buffer
x1138 gnd WL1009 net1010 vcc buffer
x1139 gnd WL1010 net1011 vcc buffer
x1140 gnd WL1011 net1012 vcc buffer
x1141 gnd WL1012 net1013 vcc buffer
x1142 gnd WL1013 net1014 vcc buffer
x1143 gnd WL1014 net1015 vcc buffer
x1144 gnd WL1015 net1016 vcc buffer
x1145 gnd WL1016 net1017 vcc buffer
x1146 gnd WL1017 net1018 vcc buffer
x1147 gnd WL1018 net1019 vcc buffer
x1148 gnd WL1019 net1020 vcc buffer
x1149 gnd WL1020 net1021 vcc buffer
x1150 gnd WL1021 net1022 vcc buffer
x1151 gnd WL1022 net1023 vcc buffer
x1152 gnd WL1023 net1024 vcc buffer
x2 vcc_bl0 PRE Blb0 Bl0 Precharge_circuit
x43 vcc_bl1 PRE Blb1 Bl1 Precharge_circuit
x44 vcc_bl2 PRE Blb2 Bl2 Precharge_circuit
x45 vcc_bl3 PRE Blb3 Bl3 Precharge_circuit
x54 vcc_bl4 PRE Blb4 Bl4 Precharge_circuit
x55 vcc_bl5 PRE Blb5 Bl5 Precharge_circuit
x56 vcc_bl6 PRE Blb6 Bl6 Precharge_circuit
x57 vcc_bl7 PRE Blb7 Bl7 Precharge_circuit
x58 vcc_bl8 PRE Blb8 Bl8 Precharge_circuit
x59 vcc_bl9 PRE Blb9 Bl9 Precharge_circuit
x60 vcc_bl10 PRE Blb10 Bl10 Precharge_circuit
x61 vcc_bl11 PRE Blb11 Bl11 Precharge_circuit
x62 vcc_bl12 PRE Blb12 Bl12 Precharge_circuit
x63 vcc_bl13 PRE Blb13 Bl13 Precharge_circuit
x72 vcc_bl14 PRE Blb14 Bl14 Precharge_circuit
x73 vcc_bl15 PRE Blb15 Bl15 Precharge_circuit
x74 vcc_bl16 PRE Blb16 Bl16 Precharge_circuit
x75 vcc_bl17 PRE Blb17 Bl17 Precharge_circuit
x76 vcc_bl18 PRE Blb18 Bl18 Precharge_circuit
x77 vcc_bl19 PRE Blb19 Bl19 Precharge_circuit
x78 vcc_bl20 PRE Blb20 Bl20 Precharge_circuit
x79 vcc_bl21 PRE Blb21 B21 Precharge_circuit
x80 vcc_bl22 PRE Blb22 Bl22 Precharge_circuit
x81 vcc_bl23 PRE Blb23 Bl23 Precharge_circuit
x82 vcc_bl24 PRE Blb24 Bl24 Precharge_circuit
x83 vcc_bl25 PRE Blb25 Bl25 Precharge_circuit
x84 vcc_bl26 PRE Blb26 Bl26 Precharge_circuit
x85 vcc_bl27 PRE Blb27 Bl27 Precharge_circuit
x86 vcc_bl28 PRE Blb28 Bl28 Precharge_circuit
x87 vcc_bl29 PRE Blb29 Bl29 Precharge_circuit
x88 vcc_bl30 PRE Blb30 Bl30 Precharge_circuit
x89 vcc_bl31 PRE Blb31 Bl31 Precharge_circuit
x1 Bl0 Blb0 writeen vcc_bl0 DataIn0 gnd_bl0 gnd write
x3 Bl1 Blb1 writeen vcc_bl1 DataIn1 gnd_bl1 gnd write
x4 Bl2 Blb2 writeen vcc_bl2 DataIn2 gnd_bl2 gnd write
x6 Bl3 Blb3 writeen vcc_bl3 DataIn3 gnd_bl3 gnd write
x7 Bl4 Blb4 writeen vcc_bl4 DataIn4 gnd_bl4 gnd write
x8 Bl5 Blb5 writeen vcc_bl5 DataIn5 gnd_bl5 gnd write
x9 Bl6 Blb6 writeen vcc_bl6 DataIn6 gnd_bl6 gnd write
x10 Bl7 Blb7 writeen vcc_bl7 DataIn7 gnd_bl7 gnd write
x11 Bl8 Blb8 writeen vcc_bl8 DataIn8 gnd_bl8 gnd write
x12 Bl9 Blb9 writeen vcc_bl9 DataIn9 gnd_bl9 gnd write
x13 Bl10 Blb10 writeen vcc_bl10 DataIn10 gnd_bl10 gnd write
x14 Bl11 Blb11 writeen vcc_bl11 DataIn11 gnd_bl11 gnd write
x15 Bl12 Blb12 writeen vcc_bl12 DataIn12 gnd_bl12 gnd write
x16 Bl13 Blb13 writeen vcc_bl13 DataIn13 gnd_bl13 gnd write
x17 Bl14 Blb14 writeen vcc_bl14 DataIn14 gnd_bl14 gnd write
x18 Bl15 Blb15 writeen vcc_bl15 DataIn15 gnd_bl15 gnd write
x19 Bl16 Blb16 writeen vcc_bl16 DataIn16 gnd_bl16 gnd write
x20 Bl17 Blb17 writeen vcc_bl17 DataIn17 gnd_bl17 gnd write
x21 Bl18 Blb18 writeen vcc_bl18 DataIn18 gnd_bl18 gnd write
x30 Bl19 Blb19 writeen vcc_bl19 DataIn19 gnd_bl19 gnd write
x31 Bl20 Blb20 writeen vcc_bl20 DataIn20 gnd_bl20 gnd write
x32 B21 Blb21 writeen vcc_bl21 DataIn21 gnd_bl21 gnd write
x33 Bl22 Blb22 writeen vcc_bl22 DataIn22 gnd_bl22 gnd write
x34 Bl23 Blb23 writeen vcc_bl23 DataIn23 gnd_bl23 gnd write
x35 Bl24 Blb24 writeen vcc_bl24 DataIn24 gnd_bl24 gnd write
x36 Bl25 Blb25 writeen vcc_bl25 DataIn25 gnd_bl25 gnd write
x37 Bl26 Blb26 writeen vcc_bl26 DataIn26 gnd_bl26 gnd write
x38 Bl27 Blb27 writeen vcc_bl27 DataIn27 gnd_bl27 gnd write
x39 Bl28 Blb28 writeen vcc_bl28 DataIn28 gnd_bl28 gnd write
x40 Bl29 Blb29 writeen vcc_bl29 DataIn29 gnd_bl29 gnd write
x41 Bl30 Blb30 writeen vcc_bl30 DataIn30 gnd_bl30 gnd write
x42 Bl31 Blb31 writeen vcc_bl31 DataIn31 gnd_bl31 gnd write
x22 vcc_bl0 DataOut0 Bl0 Blb0 readen gnd_bl0 gnd nnnsense_amp
x23 vcc_bl1 DataOut1 Bl1 Blb1 readen gnd_bl1 gnd nnnsense_amp
x24 vcc_bl2 DataOut2 Bl2 Blb2 readen gnd_bl2 gnd nnnsense_amp
x25 vcc_bl3 DataOut3 Bl3 Blb3 readen gnd_bl3 gnd nnnsense_amp
x26 vcc_bl4 DataOut4 Bl4 Blb4 readen gnd_bl4 gnd nnnsense_amp
x27 vcc_bl5 DataOut5 Bl5 Blb5 readen gnd_bl5 gnd nnnsense_amp
x28 vcc_bl6 DataOut6 Bl6 Blb6 readen gnd_bl6 gnd nnnsense_amp
x29 vcc_bl7 DataOut7 Bl7 Blb7 readen gnd_bl7 gnd nnnsense_amp
x46 vcc_bl8 DataOut8 Bl8 Blb8 readen gnd_bl8 gnd nnnsense_amp
x47 vcc_bl9 DataOut9 Bl9 Blb9 readen gnd_bl9 gnd nnnsense_amp
x48 vcc_bl10 DataOut10 Bl10 Blb10 readen gnd_bl10 gnd nnnsense_amp
x49 vcc_bl11 DataOut11 Bl11 Blb11 readen gnd_bl11 gnd nnnsense_amp
x50 vcc_bl12 DataOut12 Bl12 Blb12 readen gnd_bl12 gnd nnnsense_amp
x51 vcc_bl13 DataOut13 Bl13 Blb13 readen gnd_bl13 gnd nnnsense_amp
x52 vcc_bl14 DataOut14 Bl14 Blb14 readen gnd_bl14 gnd nnnsense_amp
x53 vcc_bl15 DataOut15 Bl15 Blb15 readen gnd_bl15 gnd nnnsense_amp
x64 vcc_bl16 DataOut16 Bl16 Blb16 readen gnd_bl16 gnd nnnsense_amp
x65 vcc_bl17 DataOut17 Bl17 Blb17 readen gnd_bl17 gnd nnnsense_amp
x66 vcc_bl18 DataOut18 Bl18 Blb18 readen gnd_bl18 gnd nnnsense_amp
x67 vcc_bl19 DataOut19 Bl19 Blb19 readen gnd_bl19 gnd nnnsense_amp
x68 vcc_bl20 DataOut20 Bl20 Blb20 readen gnd_bl20 gnd nnnsense_amp
x69 vcc_bl21 DataOut21 B21 Blb21 readen gnd_bl21 gnd nnnsense_amp
x70 vcc_bl22 DataOut22 Bl22 Blb22 readen gnd_bl22 gnd nnnsense_amp
x71 vcc_bl23 DataOut23 Bl23 Blb23 readen gnd_bl23 gnd nnnsense_amp
x90 vcc_bl24 DataOut24 Bl24 Blb24 readen gnd_bl24 gnd nnnsense_amp
x91 vcc_bl25 DataOut25 Bl25 Blb25 readen gnd_bl25 gnd nnnsense_amp
x92 vcc_bl26 DataOut26 Bl26 Blb26 readen gnd_bl26 gnd nnnsense_amp
x93 vcc_bl27 DataOut27 Bl27 Blb27 readen gnd_bl27 gnd nnnsense_amp
x94 vcc_bl28 DataOut28 Bl28 Blb28 readen gnd_bl28 gnd nnnsense_amp
x95 vcc_bl29 DataOut29 Bl29 Blb29 readen gnd_bl29 gnd nnnsense_amp
x96 vcc_bl30 DataOut30 Bl30 Blb30 readen gnd_bl30 gnd nnnsense_amp
x97 vcc_bl31 DataOut31 Bl31 Blb31 readen gnd_bl31 gnd nnnsense_amp
.ends


* expanding   symbol:
*+  /home/impact/Documents/truncation_SRAM/schematic/1bytetruncationmanagerwithand.sym # of pins=45
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/1bytetruncationmanagerwithand.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/1bytetruncationmanagerwithand.sch
.subckt 1bytetruncationmanagerwithand vcc_bl7 R7 vcc_bl6 R6 R5 vcc_bl5 R4 vcc_bl4 vcc_bl3 R3 R2
+ vcc_bl2 R1 vcc_bl1 vcc_bl0 R0 gnd_bl7 gnd_bl6 gnd_bl5 Trunk7 gnd_bl4 Trunk6 gnd_bl3 gnd_bl2 Trunk5 Trunk4
+ gnd_bl1 gnd_bl0 Trunk3 Trunk2 dataout7 Trunk1 dataout6 Trunk0 dataout5 dataout4 dataout3 dataout2 dataout1
+ Byte_Mode_EnableBar dataout0 Byte_Tail_Out Tail_In vssd1 vccd1
*.PININFO Byte_Tail_Out:O Byte_Mode_EnableBar:I R3:I R2:I R1:I R0:I R7:I R6:I R5:I R4:I Trunk3:I
*+ Trunk2:I Trunk1:I Trunk7:I Trunk6:I Trunk5:I Trunk4:I Trunk0:I dataout7:O dataout6:O dataout5:O dataout4:O
*+ gnd_bl4:B vcc_bl4:B gnd_bl5:B vcc_bl5:B gnd_bl6:B vcc_bl6:B gnd_bl7:B vcc_bl7:B gnd_bl0:B vcc_bl0:B gnd_bl1:B
*+ vcc_bl1:B gnd_bl2:B vcc_bl2:B gnd_bl3:B vcc_bl3:B dataout3:O dataout2:O dataout1:O dataout0:O Tail_In:I
*+ vssd1:B vccd1:B
x10 vccd1 Byte_Mode_EnableBar Byte_Tail_Out net1 vssd1 andun
x1 R7 R6 R5 R3 R4 R2 R1 R0 vcc_bl6 vcc_bl7 gnd_bl6 vcc_bl5 gnd_bl7 vcc_bl3 vcc_bl4 Tail_In gnd_bl5
+ gnd_bl4 gnd_bl3 dataout6 dataout7 dataout5 dataout4 dataout3 vccd1 vssd1 vcc_bl2 gnd_bl2 dataout2 Trunk7
+ Trunk6 Trunk5 Trunk4 vcc_bl1 Trunk3 gnd_bl1 Trunk2 Trunk1 Trunk0 dataout1 vcc_bl0 gnd_bl0 net1 dataout0
+ 1byte_truncationmanager
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/32x32_truncation_sram.sym #
*+ of pins=161
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/32x32_truncation_sram.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/32x32_truncation_sram.sch
.subckt 32x32_truncation_sram vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3
+ vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10
+ gnd_bl10 vcc_bl11 gnd_bl11 vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 vcc_bl16
+ gnd_bl16 vcc_bl17 gnd_bl17 vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20 vcc_bl21 gnd_bl21 vcc_bl22
+ gnd_bl22 vcc_bl23 gnd_bl23 vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26 vcc_bl27 gnd_bl27 vcc_bl28
+ gnd_bl28 vcc_bl29 gnd_bl29 vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 Wl0 Wl1 Wl2 Wl3 Wl4 Wl5 Wl6 Wl7 Wl8 Wl9 Wl10
+ Wl11 Wl12 Wl13 Wl14 Wl15 Wl16 Wl17 Wl18 Wl19 Wl20 Wl21 Wl22 Wl23 Wl24 Wl25 Wl26 Wl27 Wl28 Wl29 Wl30 Wl31
+ Blb13 Bl13 Blb12 Blb11 Bl11 Blb10 Blb9 Bl9 Blb8 Bl8 Blb31 Bl31 Blb30 Blb7 Bl7 Blb6 Bl6 Blb28 Blb5 Bl10
+ Blb27 Blb26 Bl5 Bl12 Blb4 Bl4 Blb24 Bl14 Blb3 Blb23 Bl23 Blb22 Bl3 Blb2 Blb21 Blb20 Bl2 Bl20 Blb19 Bl19
+ Blb18 Bl21 Blb1 Bl22 Bl18 Blb17 Bl17 Bl24 Blb16 Bl25 Blb25 Bl26 Bl16 Bl27 Blb15 Bl28 Bl15 Bl29 Blb29 Bl30
+ Blb14 Bl1 Blb0 Bl0 gnd
*.PININFO Wl0:I Wl1:I Wl2:I Wl3:I Wl4:I Wl5:I Wl6:I Wl7:I Wl8:I Wl9:I Wl10:I Wl11:I Wl12:I Wl13:I
*+ Wl14:I Wl15:I Wl16:I Wl17:I Wl18:I Wl19:I Wl20:I Wl21:I Wl22:I Wl23:I Wl24:I Wl25:I Wl26:I Wl27:I Wl28:I
*+ Wl29:I Wl30:I Wl31:I Bl0:B Blb0:B Bl1:B Blb1:B Bl2:B Blb2:B Bl3:B Blb3:B Bl4:B Blb4:B Bl5:B Blb5:B Bl6:B
*+ Blb6:B Bl7:B Blb7:B Bl8:B Blb8:B Bl9:B Blb9:B Bl10:B Blb10:B Bl11:B Blb11:B Bl12:B Blb12:B Bl13:B Blb13:B
*+ Bl14:B Blb14:B Bl15:B Blb15:B Bl16:B Blb16:B Bl17:B Blb17:B Bl18:B Blb18:B Bl19:B Blb19:B Bl20:B Blb20:B
*+ Bl21:B Blb21:B Bl22:B Blb22:B Bl23:B Blb23:B Bl24:B Blb24:B Bl25:B Blb25:B Bl26:B Blb26:B Bl27:B Blb27:B
*+ Bl28:B Blb28:B Bl29:B Blb29:B Bl30:B Blb30:B Bl31:B Blb31:B vcc_bl0:B vcc_bl1:B vcc_bl2:B vcc_bl3:B
*+ gnd_bl0:B gnd_bl1:B gnd_bl2:B gnd_bl3:B vcc_bl4:B vcc_bl5:B vcc_bl6:B vcc_bl7:B gnd_bl4:B gnd_bl5:B gnd_bl6:B
*+ gnd_bl7:B vcc_bl8:B vcc_bl9:B vcc_bl10:B vcc_bl11:B gnd_bl8:B gnd_bl9:B gnd_bl10:B gnd_bl11:B vcc_bl12:B
*+ vcc_bl13:B vcc_bl14:B vcc_bl15:B gnd_bl12:B gnd_bl13:B gnd_bl14:B gnd_bl15:B vcc_bl16:B vcc_bl17:B vcc_bl18:B
*+ vcc_bl19:B gnd_bl16:B gnd_bl17:B gnd_bl18:B gnd_bl19:B vcc_bl20:B vcc_bl21:B vcc_bl22:B vcc_bl23:B gnd_bl20:B
*+ gnd_bl21:B gnd_bl22:B gnd_bl23:B vcc_bl24:B vcc_bl25:B vcc_bl26:B vcc_bl27:B gnd_bl24:B gnd_bl25:B gnd_bl26:B
*+ gnd_bl27:B vcc_bl28:B vcc_bl29:B vcc_bl30:B vcc_bl31:B gnd_bl28:B gnd_bl29:B gnd_bl30:B gnd_bl31:B gnd:B
x1 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 Wl0 Wl1 Wl2 Wl3 Wl4 Wl5 Wl6 Wl7 Wl8
+ Wl9 Wl10 Wl11 Wl12 Wl13 Wl14 Wl15 Blb5 Bl5 Blb4 Blb3 Blb15 Bl15 Blb14 Bl4 Bl3 Blb2 Bl2 Bl6 Blb12 Blb1
+ Blb11 Bl11 Blb10 Bl1 Bl10 Blb9 Bl9 Blb8 Bl8 Bl12 Blb7 Bl13 Blb13 Bl14 Bl7 Blb6 Blb0 Bl0 gnd 16x16_sram
x2 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17 vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20
+ vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23 vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26
+ vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29 vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 Wl0 Wl1 Wl2 Wl3
+ Wl4 Wl5 Wl6 Wl7 Wl8 Wl9 Wl10 Wl11 Wl12 Wl13 Wl14 Wl15 Blb21 Bl21 Blb20 Blb19 Blb31 Bl31 Blb30 Bl20 Bl19
+ Blb18 Bl18 Bl22 Blb28 Blb17 Blb27 Bl27 Blb26 Bl17 Bl26 Blb25 Bl25 Blb24 Bl24 Bl28 Blb23 Bl29 Blb29 Bl30
+ Bl23 Blb22 Blb16 Bl16 gnd 16x16_sram
x3 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11
+ vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 Wl16 Wl17 Wl18 Wl19 Wl20 Wl21 Wl22
+ Wl23 Wl24 Wl25 Wl26 Wl27 Wl28 Wl29 Wl30 Wl31 Blb5 Bl5 Blb4 Blb3 Blb15 Bl15 Blb14 Bl4 Bl3 Blb2 Bl2 Bl6
+ Blb12 Blb1 Blb11 Bl11 Blb10 Bl1 Bl10 Blb9 Bl9 Blb8 Bl8 Bl12 Blb7 Bl13 Blb13 Bl14 Bl7 Blb6 Blb0 Bl0 gnd
+ 16x16_sram
x4 vcc_bl16 gnd_bl16 vcc_bl17 gnd_bl17 vcc_bl18 gnd_bl18 vcc_bl19 gnd_bl19 vcc_bl20 gnd_bl20
+ vcc_bl21 gnd_bl21 vcc_bl22 gnd_bl22 vcc_bl23 gnd_bl23 vcc_bl24 gnd_bl24 vcc_bl25 gnd_bl25 vcc_bl26 gnd_bl26
+ vcc_bl27 gnd_bl27 vcc_bl28 gnd_bl28 vcc_bl29 gnd_bl29 vcc_bl30 gnd_bl30 vcc_bl31 gnd_bl31 Wl16 Wl17 Wl18
+ Wl19 Wl20 Wl21 Wl22 Wl23 Wl24 Wl25 Wl26 Wl27 Wl28 Wl29 Wl30 Wl31 Blb21 Bl21 Blb20 Blb19 Blb31 Bl31 Blb30
+ Bl20 Bl19 Blb18 Bl18 Bl22 Blb28 Blb17 Blb27 Bl27 Blb26 Bl17 Bl26 Blb25 Bl25 Blb24 Bl24 Bl28 Blb23 Bl29
+ Blb29 Bl30 Bl23 Blb22 Blb16 Bl16 gnd 16x16_sram
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/buffer.sym # of pins=4
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/buffer.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/buffer.sch
.subckt buffer gnd In Out vcc
*.PININFO In:B Out:B gnd:B vcc:B
XM6 Out net1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM1 net1 In gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM10 Out net1 vcc vcc sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM5 net1 In vcc vcc sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/Precharge_circuit.sym # of
*+ pins=4
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/Precharge_circuit.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/Precharge_circuit.sch
.subckt Precharge_circuit vcc PreB Blb Bl
*.PININFO vcc:B PreB:I Bl:B Blb:B
XM9 Blb PreB vcc vcc sky130_fd_pr__pfet_01v8 L=0.18 W=0.72 nf=1 m=1
XM10 Bl PreB vcc vcc sky130_fd_pr__pfet_01v8 L=0.18 W=0.72 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/write.sym # of pins=7
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/write.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/write.sch
.subckt write Bl Blb Wen vdd DATA gnd_virtual gnd
*.PININFO vdd:B gnd:B Bl:B Blb:B Wen:B DATA:B gnd_virtual:B
XM7 Bl_X Wen Bl gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM1 Blb Wen Blb_X gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
x1 vdd Blb_X Bl_X gnd gnd_virtual inverter_virtual
x2 vdd Inv_X DATA gnd gnd_virtual inverter_virtual
x3 vdd Bl_X Inv_X gnd gnd_virtual inverter_virtual
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/nnnsense_amp.sym # of pins=7
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/nnnsense_amp.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/nnnsense_amp.sch
.subckt nnnsense_amp vdd BlOut Bl Blb readEn gnd_virtual gnd
*.PININFO vdd:B gnd:B readEn:B Blb:B Bl:B BlOut:B gnd_virtual:B
XM1 net3 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=0.84 nf=1 m=1
XM2 net3 Bl net2 gnd sky130_fd_pr__nfet_01v8 L=0.18 W=0.42 nf=1 m=1
XM3 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=0.84 nf=1 m=1
XM4 net1 Blb net2 gnd sky130_fd_pr__nfet_01v8 L=0.18 W=0.42 nf=1 m=1
XM5 BlOut net3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=0.84 nf=1 m=1
XM6 BlOut net3 gnd_virtual gnd sky130_fd_pr__nfet_01v8 L=0.18 W=0.42 nf=1 m=1
XM7 net2 readEn gnd_virtual gnd sky130_fd_pr__nfet_01v8 L=0.18 W=1.26 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/andun.sym # of pins=5
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/andun.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/andun.sch
.subckt andun vccd1 A Out B vssd1
*.PININFO Out:O A:I B:I vssd1:B vccd1:B
x1 vccd1 net1 A B vssd1 nandAB
x2 vccd1 net1 Out vssd1 inverter_symbol
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/1byte_truncationmanager.sym
*+ # of pins=44
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/1byte_truncationmanager.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/1byte_truncationmanager.sch
.subckt 1byte_truncationmanager R7 R6 R5 R3 R4 R2 R1 R0 vcc_bl6 vcc_bl7 gnd_bl6 vcc_bl5 gnd_bl7
+ vcc_bl3 vcc_bl4 Tail_In gnd_bl5 gnd_bl4 gnd_bl3 dataout6 dataout7 dataout5 dataout4 dataout3 vccd1 vssd1
+ vcc_bl2 gnd_bl2 dataout2 Trunk7 Trunk6 Trunk5 Trunk4 vcc_bl1 Trunk3 gnd_bl1 Trunk2 Trunk1 Trunk0 dataout1
+ vcc_bl0 gnd_bl0 Tail_Out dataout0
*.PININFO vcc_bl0:B gnd_bl0:B vcc_bl1:B gnd_bl1:B vcc_bl2:B gnd_bl2:B vcc_bl3:B gnd_bl3:B dataout3:O
*+ dataout2:O dataout1:O Trunk3:I Trunk2:I Trunk1:I Trunk0:I R3:I R2:I R1:I R0:I Tail_In:I R4:I R5:I R6:I R7:I
*+ vcc_bl4:B gnd_bl4:B vcc_bl5:B gnd_bl5:B vcc_bl6:B gnd_bl6:B vcc_bl7:B gnd_bl7:B dataout7:O dataout6:O
*+ dataout5:O dataout4:O Trunk7:I Trunk6:I Trunk5:I Trunk4:I Tail_Out:O vccd1:B vssd1:B dataout0:O
x1 Trunk7 vcc_bl7 gnd_bl7 Tail_In net7 vccd1 vssd1 R7 dataout7 truncation_manager
x2 Trunk6 vcc_bl6 gnd_bl6 net7 net6 vccd1 vssd1 R6 dataout6 truncation_manager
x3 Trunk5 vcc_bl5 gnd_bl5 net6 net5 vccd1 vssd1 R5 dataout5 truncation_manager
x4 Trunk4 vcc_bl4 gnd_bl4 net5 net4 vccd1 vssd1 R4 dataout4 truncation_manager
x5 Trunk3 vcc_bl3 gnd_bl3 net4 net1 vccd1 vssd1 R3 dataout3 truncation_manager
x6 Trunk2 vcc_bl2 gnd_bl2 net1 net2 vccd1 vssd1 R2 dataout2 truncation_manager
x7 Trunk1 vcc_bl1 gnd_bl1 net2 net3 vccd1 vssd1 R1 dataout1 truncation_manager
x8 Trunk0 vcc_bl0 gnd_bl0 net3 Tail_Out vccd1 vssd1 R0 dataout0 truncation_manager
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/16x16_sram.sym # of pins=81
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/16x16_sram.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/16x16_sram.sch
.subckt 16x16_sram vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4
+ vcc_bl5 gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11
+ gnd_bl11 vcc_bl12 gnd_bl12 vcc_bl13 gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 Wl0 Wl1 Wl2 Wl3 Wl4 Wl5 Wl6
+ Wl7 Wl8 Wl9 Wl10 Wl11 Wl12 Wl13 Wl14 Wl15 Blb5 Bl5 Blb4 Blb3 Blb15 Bl15 Blb14 Bl4 Bl3 Blb2 Bl2 Bl6
+ Blb12 Blb1 Blb11 Bl11 Blb10 Bl1 Bl10 Blb9 Bl9 Blb8 Bl8 Bl12 Blb7 Bl13 Blb13 Bl14 Bl7 Blb6 Blb0 Bl0 gnd
*.PININFO Wl0:I Wl1:I Wl2:I Wl3:I Wl4:I Wl5:I Wl6:I Wl7:I Wl8:I Wl9:I Wl10:I Wl11:I Wl12:I Wl13:I
*+ Wl14:I Wl15:I Bl0:B Blb0:B Bl1:B Blb1:B Bl2:B Blb2:B Bl3:B Blb3:B Bl4:B Blb4:B Bl5:B Blb5:B Bl6:B Blb6:B
*+ Bl7:B Blb7:B Bl8:B Blb8:B Bl9:B Blb9:B Bl10:B Blb10:B Bl11:B Blb11:B Bl12:B Blb12:B Bl13:B Blb13:B Bl14:B
*+ Blb14:B Bl15:B Blb15:B vcc_bl0:B vcc_bl1:B vcc_bl2:B vcc_bl3:B gnd_bl0:B gnd_bl1:B gnd_bl2:B gnd_bl3:B
*+ vcc_bl4:B vcc_bl5:B vcc_bl6:B vcc_bl7:B gnd_bl4:B gnd_bl5:B gnd_bl6:B gnd_bl7:B vcc_bl8:B vcc_bl9:B
*+ vcc_bl10:B vcc_bl11:B gnd_bl8:B gnd_bl9:B gnd_bl10:B gnd_bl11:B vcc_bl12:B vcc_bl13:B vcc_bl14:B vcc_bl15:B
*+ gnd_bl12:B gnd_bl13:B gnd_bl14:B gnd_bl15:B gnd:B
x1 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 Bl3 Blb2 Bl2 Blb7 Blb1 Bl7 Blb6 Bl1 Bl6 Blb5 Blb0 Bl5 Blb4 Bl0 Bl4 Blb3 Wl0
+ Wl1 Wl2 Wl3 Wl4 Wl5 Wl6 Wl7 gnd 8x8_truncation_sram
x2 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11 vcc_bl12 gnd_bl12 vcc_bl13
+ gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 Bl11 Blb10 Bl10 Blb15 Blb9 Bl15 Blb14 Bl9 Bl14 Blb13 Blb8 Bl13
+ Blb12 Bl8 Bl12 Blb11 Wl0 Wl1 Wl2 Wl3 Wl4 Wl5 Wl6 Wl7 gnd 8x8_truncation_sram
x3 vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4 gnd_bl4 vcc_bl5 gnd_bl5
+ vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 Bl3 Blb2 Bl2 Blb7 Blb1 Bl7 Blb6 Bl1 Bl6 Blb5 Blb0 Bl5 Blb4 Bl0 Bl4 Blb3 Wl8
+ Wl9 Wl10 Wl11 Wl12 Wl13 Wl14 Wl15 gnd 8x8_truncation_sram
x4 vcc_bl8 gnd_bl8 vcc_bl9 gnd_bl9 vcc_bl10 gnd_bl10 vcc_bl11 gnd_bl11 vcc_bl12 gnd_bl12 vcc_bl13
+ gnd_bl13 vcc_bl14 gnd_bl14 vcc_bl15 gnd_bl15 Bl11 Blb10 Bl10 Blb15 Blb9 Bl15 Blb14 Bl9 Bl14 Blb13 Blb8 Bl13
+ Blb12 Bl8 Bl12 Blb11 Wl8 Wl9 Wl10 Wl11 Wl12 Wl13 Wl14 Wl15 gnd 8x8_truncation_sram
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/inverter_virtual.sym # of
*+ pins=5
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/inverter_virtual.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/inverter_virtual.sch
.subckt inverter_virtual vccd1 Out In vssd1 gnd_virtual
*.PININFO vccd1:B vssd1:B gnd_virtual:B Out:B In:B
XM8 Out In vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM9 Out In gnd_virtual vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/nandAB.sym # of pins=5
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/nandAB.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/nandAB.sch
.subckt nandAB vccd1 Out A B vssd1
*.PININFO Out:O A:I vccd1:B vssd1:B B:I
XM1 Out B vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=.84 nf=1 m=1
XM2 Out A vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=.84 nf=1 m=1
XM6 net1 B vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM9 Out A net1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/inverter_symbol.sym # of
*+ pins=4
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/inverter_symbol.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/inverter_symbol.sch
.subckt inverter_symbol vccd1 In Out vssd1
*.PININFO In:I Out:O vccd1:B vssd1:B
XM3 Out In vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM4 Out In vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/truncation_manager.sym # of
*+ pins=9
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/truncation_manager.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/truncation_manager.sch
.subckt truncation_manager Head vcc_Bl gnd_Bl Tail_In Tail_Out vccd1 vssd1 Bl ReadOut
*.PININFO vccd1:B Head:I Bl:I Tail_In:I Tail_Out:O gnd_Bl:B vcc_Bl:B vssd1:B ReadOut:O
x2 vccd1 Tail_Out vcc_Bl gnd_Bl vssd1 final_power_gate
x1 vssd1 vccd1 net1 Head Tail_Out Tail_In schem_truncationunit
x3 vccd1 net1 Tail_Out ReadOut Bl vssd1 mysch_mux
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/8x8_truncation_sram.sym # of
*+ pins=41
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/8x8_truncation_sram.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/8x8_truncation_sram.sch
.subckt 8x8_truncation_sram vcc_bl0 gnd_bl0 vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 vcc_bl4
+ gnd_bl4 vcc_bl5 gnd_bl5 vcc_bl6 gnd_bl6 vcc_bl7 gnd_bl7 Bl3 Blb2 Bl2 Blb7 Blb1 Bl7 Blb6 Bl1 Bl6 Blb5 Blb0
+ Bl5 Blb4 Bl0 Bl4 Blb3 Wl0 Wl1 Wl2 Wl3 Wl4 Wl5 Wl6 Wl7 gnd
*.PININFO Wl0:I Wl1:I Wl2:I Wl7:I Wl3:I Wl4:I Wl5:I Wl6:I Bl0:B Blb0:B Bl1:B Blb1:B Bl2:B Blb2:B
*+ Bl3:B Blb3:B Bl4:B Blb4:B Bl5:B Blb5:B Bl6:B Blb6:B Bl7:B Blb7:B vcc_bl0:B vcc_bl1:B vcc_bl2:B vcc_bl3:B
*+ gnd_bl0:B gnd_bl1:B gnd_bl2:B gnd_bl3:B vcc_bl4:B vcc_bl5:B vcc_bl6:B vcc_bl7:B gnd_bl4:B gnd_bl5:B gnd_bl6:B
*+ gnd_bl7:B gnd:B
x1 vcc_bl0 gnd_bl0 Bl1 Blb3 Blb0 Bl3 Blb2 Bl0 Bl2 Blb1 Wl0 Wl1 Wl2 Wl3 vcc_bl1 gnd_bl1 vcc_bl2
+ gnd_bl2 vcc_bl3 gnd_bl3 gnd 4x4_truncation_sram
x2 vcc_bl4 gnd_bl4 Bl5 Blb7 Blb4 Bl7 Blb6 Bl4 Bl6 Blb5 Wl0 Wl1 Wl2 Wl3 vcc_bl5 gnd_bl5 vcc_bl6
+ gnd_bl6 vcc_bl7 gnd_bl7 gnd 4x4_truncation_sram
x3 vcc_bl0 gnd_bl0 Bl1 Blb3 Blb0 Bl3 Blb2 Bl0 Bl2 Blb1 Wl4 Wl5 Wl6 Wl7 vcc_bl1 gnd_bl1 vcc_bl2
+ gnd_bl2 vcc_bl3 gnd_bl3 gnd 4x4_truncation_sram
x4 vcc_bl4 gnd_bl4 Bl5 Blb7 Blb4 Bl7 Blb6 Bl4 Bl6 Blb5 Wl4 Wl5 Wl6 Wl7 vcc_bl5 gnd_bl5 vcc_bl6
+ gnd_bl6 vcc_bl7 gnd_bl7 gnd 4x4_truncation_sram
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/final_power_gate.sym # of
*+ pins=5
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/final_power_gate.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/final_power_gate.sch
.subckt final_power_gate vcc enb vcc_out gnd_out gnd
*.PININFO enb:I vcc:B gnd:B vcc_out:B gnd_out:B
XM5 net1 enb gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net1 enb vcc vcc sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 vcc_out enb vcc vcc sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=8 m=1
XM2 gnd_out net1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=8 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/schem_truncationunit.sym #
*+ of pins=6
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/schem_truncationunit.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/schem_truncationunit.sch
.subckt schem_truncationunit gnd vcc Bl head tail_signal tail
*.PININFO head:I tail:I tail_signal:O gnd:B Bl:O vcc:B
XM1 Bl net2 net1 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
x4 vcc head net3 gnd inverter_symbol
x1 vcc net1 tail net3 gnd nandAB
x2 vcc tail_signal head tail gnd or_gate
x3 vcc net2 tail head gnd or_gate
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/mysch_mux.sym # of pins=6
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/mysch_mux.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/mysch_mux.sch
.subckt mysch_mux vccd1 A1 S X A0 vssd1
*.PININFO vccd1:B A1:I X:O vssd1:B S:I A0:I
x1 vccd1 S net3 A1 vssd1 andun
x3 vccd1 X net3 net2 vssd1 or_gate
x4 vccd1 A0 net2 net1 vssd1 andun
x2 vccd1 S net1 vssd1 inverter_symbol
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/4x4_truncation_sram.sym # of
*+ pins=21
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/4x4_truncation_sram.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/4x4_truncation_sram.sch
.subckt 4x4_truncation_sram vcc_bl0 gnd_bl0 bl1 blb3 blb0 bl3 blb2 bl0 bl2 blb1 Wl0 Wl1 Wl2 Wl3
+ vcc_bl1 gnd_bl1 vcc_bl2 gnd_bl2 vcc_bl3 gnd_bl3 gnd
*.PININFO Wl0:I Wl1:I Wl2:I Wl3:I bl0:B blb0:B bl1:B blb1:B bl2:B blb2:B bl3:B blb3:B vcc_bl0:B
*+ vcc_bl1:B vcc_bl2:B vcc_bl3:B gnd_bl0:B gnd_bl1:B gnd_bl2:B gnd_bl3:B gnd:B
x1 bl1 blb1 blb0 bl0 Wl0 Wl1 vcc_bl0 gnd_bl1 vcc_bl1 gnd_bl0 gnd 2x2_truncation_sram
x2 bl3 blb3 blb2 bl2 Wl0 Wl1 vcc_bl2 gnd_bl3 vcc_bl3 gnd_bl2 gnd 2x2_truncation_sram
x3 bl1 blb1 blb0 bl0 Wl2 Wl3 vcc_bl0 gnd_bl1 vcc_bl1 gnd_bl0 gnd 2x2_truncation_sram
x4 bl3 blb3 blb2 bl2 Wl2 Wl3 vcc_bl2 gnd_bl3 vcc_bl3 gnd_bl2 gnd 2x2_truncation_sram
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/or_gate.sym # of pins=5
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/or_gate.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/or_gate.sch
.subckt or_gate vccd1 Out A B vssd1
*.PININFO Out:O A:I vccd1:B vssd1:B B:I
XM1 net1 A vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=.84 nf=1 m=1
XM2 net2 B net1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=.84 nf=1 m=1
XM9 net2 B vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM3 net2 A vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM6 Out net2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM7 Out net2 vccd1 vccd1 sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/2x2_truncation_sram.sym # of
*+ pins=11
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/2x2_truncation_sram.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/2x2_truncation_sram.sch
.subckt 2x2_truncation_sram Bl1 Blb1 Blb0 Bl0 Wl0 Wl1 vcc_Bl0 gnd_Bl1 vcc_Bl1 gnd_Bl0 gnd
*.PININFO Blb0:B Bl0:B Blb1:B Bl1:B Wl0:I Wl1:I gnd_Bl0:B vcc_Bl0:B vcc_Bl1:B gnd_Bl1:B gnd:B
x1 Wl0 vcc_Bl0 Blb0 Bl0 gnd_Bl0 gnd 6t_sram_virtual
x2 Wl0 vcc_Bl1 Blb1 Bl1 gnd_Bl1 gnd 6t_sram_virtual
x3 Wl1 vcc_Bl0 Blb0 Bl0 gnd_Bl0 gnd 6t_sram_virtual
x4 Wl1 vcc_Bl1 Blb1 Bl1 gnd_Bl1 gnd 6t_sram_virtual
.ends


* expanding   symbol:  /home/impact/Documents/truncation_SRAM/schematic/6t_sram_virtual.sym # of
*+ pins=6
** sym_path: /home/impact/Documents/truncation_SRAM/schematic/6t_sram_virtual.sym
** sch_path: /home/impact/Documents/truncation_SRAM/schematic/6t_sram_virtual.sch
.subckt 6t_sram_virtual Wl vcc_virtual Blb Bl gnd_virtual gnd
*.PININFO gnd_virtual:B vcc_virtual:B Blb:B Bl:B Wl:I gnd:B
XM1 Qb Q vcc_virtual vcc_virtual sky130_fd_pr__pfet_01v8 L=0.15 W=0.55 nf=1 m=1
XM2 Qb Q gnd_virtual gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=1 m=1
XM3 Q Qb vcc_virtual vcc_virtual sky130_fd_pr__pfet_01v8 L=0.15 W=0.55 nf=1 m=1
XM4 Q Qb gnd_virtual gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=1 m=1
XM7 Q Wl Bl gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 Qb Wl Blb gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends

.end
