VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO privacy_SRAM
  CLASS BLOCK ;
  FOREIGN privacy_SRAM ;
  ORIGIN -42.000 -8.150 ;
  SIZE 156.000 BY 230.000 ;
  PIN WL0
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 164.350 44.000 164.950 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 162.550 44.000 163.150 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 160.750 44.000 161.350 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 158.950 44.000 159.550 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 157.150 44.000 157.750 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 155.350 44.000 155.950 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 153.550 44.000 154.150 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 151.750 44.000 152.350 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 149.950 44.000 150.550 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 148.150 44.000 148.750 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 146.350 44.000 146.950 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 144.550 44.000 145.150 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 142.750 44.000 143.350 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 140.950 44.000 141.550 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 139.150 44.000 139.750 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 137.350 44.000 137.950 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 135.550 44.000 136.150 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 133.750 44.000 134.350 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 131.950 44.000 132.550 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 130.150 44.000 130.750 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 128.350 44.000 128.950 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 126.550 44.000 127.150 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 124.750 44.000 125.350 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 122.950 44.000 123.550 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 121.150 44.000 121.750 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 119.350 44.000 119.950 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 117.550 44.000 118.150 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 115.750 44.000 116.350 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 113.950 44.000 114.550 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 112.150 44.000 112.750 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 110.350 44.000 110.950 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 108.550 44.000 109.150 ;
    END
  END WL31
  PIN WL32
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 100.500 44.000 101.100 ;
    END
  END WL32
  PIN WL33
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 98.900 44.000 99.500 ;
    END
  END WL33
  PIN WL34
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 97.300 44.000 97.900 ;
    END
  END WL34
  PIN WL35
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 95.700 44.000 96.300 ;
    END
  END WL35
  PIN WL36
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 94.100 44.000 94.700 ;
    END
  END WL36
  PIN WL37
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 92.500 44.000 93.100 ;
    END
  END WL37
  PIN WL38
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 90.900 44.000 91.500 ;
    END
  END WL38
  PIN WL39
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 89.300 44.000 89.900 ;
    END
  END WL39
  PIN WL40
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 87.700 44.000 88.300 ;
    END
  END WL40
  PIN WL41
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 86.100 44.000 86.700 ;
    END
  END WL41
  PIN WL42
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 84.500 44.000 85.100 ;
    END
  END WL42
  PIN WL43
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 82.900 44.000 83.500 ;
    END
  END WL43
  PIN WL44
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 81.300 44.000 81.900 ;
    END
  END WL44
  PIN WL45
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 79.700 44.000 80.300 ;
    END
  END WL45
  PIN WL46
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 78.100 44.000 78.700 ;
    END
  END WL46
  PIN WL47
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 76.500 44.000 77.100 ;
    END
  END WL47
  PIN WL48
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 74.900 44.000 75.500 ;
    END
  END WL48
  PIN WL49
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 73.300 44.000 73.900 ;
    END
  END WL49
  PIN WL50
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 71.700 44.000 72.300 ;
    END
  END WL50
  PIN WL51
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 70.100 44.000 70.700 ;
    END
  END WL51
  PIN WL52
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 68.500 44.000 69.100 ;
    END
  END WL52
  PIN WL53
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 66.900 44.000 67.500 ;
    END
  END WL53
  PIN WL54
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 65.300 44.000 65.900 ;
    END
  END WL54
  PIN WL55
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 63.700 44.000 64.300 ;
    END
  END WL55
  PIN WL56
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 62.100 44.000 62.700 ;
    END
  END WL56
  PIN WL57
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 60.500 44.000 61.100 ;
    END
  END WL57
  PIN WL58
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 58.900 44.000 59.500 ;
    END
  END WL58
  PIN WL59
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 57.300 44.000 57.900 ;
    END
  END WL59
  PIN WL60
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 55.700 44.000 56.300 ;
    END
  END WL60
  PIN WL61
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 54.100 44.000 54.700 ;
    END
  END WL61
  PIN WL62
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 52.500 44.000 53.100 ;
    END
  END WL62
  PIN WL63
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 50.900 44.000 51.500 ;
    END
  END WL63
  PIN DataOut0
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 99.300 236.100 99.750 238.100 ;
    END
  END DataOut0
  PIN DataOut1
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 106.050 236.150 106.500 238.150 ;
    END
  END DataOut1
  PIN DataOut2
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 112.800 236.150 113.250 238.150 ;
    END
  END DataOut2
  PIN DataOut3
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 119.550 236.150 120.000 238.150 ;
    END
  END DataOut3
  PIN DataOut4
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 126.300 236.150 126.750 238.150 ;
    END
  END DataOut4
  PIN DataOut5
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 133.050 236.150 133.500 238.150 ;
    END
  END DataOut5
  PIN DataOut6
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 139.800 236.150 140.250 238.150 ;
    END
  END DataOut6
  PIN DataOut7
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 146.550 236.150 147.000 238.150 ;
    END
  END DataOut7
  PIN DataOut8
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 153.300 236.150 153.750 238.150 ;
    END
  END DataOut8
  PIN DataOut9
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 160.050 236.150 160.500 238.150 ;
    END
  END DataOut9
  PIN DataIn0
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 93.350 236.150 94.050 238.150 ;
    END
  END DataIn0
  PIN DataIn1
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 100.100 236.150 100.800 238.150 ;
    END
  END DataIn1
  PIN DataIn2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 106.850 236.150 107.550 238.150 ;
    END
  END DataIn2
  PIN DataIn3
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 113.600 236.150 114.300 238.150 ;
    END
  END DataIn3
  PIN DataIn4
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 120.350 236.150 121.050 238.150 ;
    END
  END DataIn4
  PIN DataIn5
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 127.100 236.150 127.800 238.150 ;
    END
  END DataIn5
  PIN DataIn6
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 133.850 236.150 134.550 238.150 ;
    END
  END DataIn6
  PIN DataIn7
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 140.600 236.150 141.300 238.150 ;
    END
  END DataIn7
  PIN DataIn8
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 147.350 236.150 148.050 238.150 ;
    END
  END DataIn8
  PIN DataIn9
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 154.100 236.150 154.800 238.150 ;
    END
  END DataIn9
  PIN write_en
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 174.100 44.000 174.700 ;
    END
  END write_en
  PIN read_en
    ANTENNAGATEAREA 2.268000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 171.450 44.000 172.050 ;
    END
  END read_en
  PIN vccd1
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 44.000 8.150 48.000 10.150 ;
        RECT 93.700 9.500 94.250 10.150 ;
        RECT 96.450 9.500 97.000 10.150 ;
        RECT 99.200 9.500 99.750 10.150 ;
        RECT 101.950 9.500 102.500 10.150 ;
        RECT 104.700 9.500 105.250 10.150 ;
        RECT 107.450 9.500 108.000 10.150 ;
        RECT 192.000 8.150 196.000 10.150 ;
      LAYER via2 ;
        RECT 44.750 8.900 47.250 10.150 ;
        RECT 93.800 9.600 94.150 10.150 ;
        RECT 96.550 9.600 96.900 10.150 ;
        RECT 99.300 9.600 99.650 10.150 ;
        RECT 102.050 9.600 102.400 10.150 ;
        RECT 104.800 9.600 105.150 10.150 ;
        RECT 107.550 9.600 107.900 10.150 ;
        RECT 192.750 8.900 195.250 10.150 ;
      LAYER met3 ;
        RECT 42.000 232.150 198.000 236.150 ;
        RECT 42.000 10.150 44.000 12.150 ;
        RECT 196.000 10.150 198.000 12.150 ;
        RECT 42.000 8.150 198.000 10.150 ;
    END
  END vccd1
  PIN vssd1
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 42.000 223.150 198.000 227.150 ;
        RECT 42.000 17.150 44.000 21.150 ;
        RECT 196.000 17.150 198.000 21.150 ;
    END
  END vssd1
  PIN vccd2
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 42.000 214.150 198.000 218.150 ;
        RECT 42.000 26.150 44.000 30.150 ;
        RECT 196.000 26.150 198.000 30.150 ;
    END
  END vccd2
  PIN vssd2
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 42.000 205.150 198.000 209.150 ;
        RECT 42.000 35.150 44.000 39.150 ;
        RECT 196.000 35.150 198.000 39.150 ;
    END
  END vssd2
  PIN PreB
    ANTENNAGATEAREA 2.592000 ;
    PORT
      LAYER met3 ;
        RECT 42.000 46.000 44.000 46.600 ;
    END
  END PreB
  OBS
      LAYER li1 ;
        RECT 80.660 44.510 160.520 200.650 ;
      LAYER met1 ;
        RECT 53.700 44.510 168.450 200.650 ;
      LAYER met2 ;
        RECT 44.000 10.150 196.000 236.150 ;
      LAYER met3 ;
        RECT 44.000 10.150 196.000 189.350 ;
  END
END privacy_SRAM
END LIBRARY

