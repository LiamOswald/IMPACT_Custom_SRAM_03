VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_IMPACT_HEAD
  CLASS BLOCK ;
  FOREIGN user_proj_IMPACT_HEAD ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 3000.000 ;
  PIN Byte_Mode_Enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1831.960 4.000 1832.560 ;
    END
  END Byte_Mode_Enable
  PIN Byte_Select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END Byte_Select[0]
  PIN Byte_Select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END Byte_Select[1]
  PIN Data_In[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END Data_In[0]
  PIN Data_In[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END Data_In[1]
  PIN Data_In[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END Data_In[2]
  PIN Data_In[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END Data_In[3]
  PIN Data_In[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 4.000 ;
    END
  END Data_In[4]
  PIN Data_In[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END Data_In[5]
  PIN Data_In[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1105.470 0.000 1105.750 4.000 ;
    END
  END Data_In[6]
  PIN Data_In[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1201.610 0.000 1201.890 4.000 ;
    END
  END Data_In[7]
  PIN Data_In_Enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END Data_In_Enable
  PIN Data_Out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END Data_Out[0]
  PIN Data_Out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1393.890 0.000 1394.170 4.000 ;
    END
  END Data_Out[1]
  PIN Data_Out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END Data_Out[2]
  PIN Data_Out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1586.170 0.000 1586.450 4.000 ;
    END
  END Data_Out[3]
  PIN Data_Out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1682.310 0.000 1682.590 4.000 ;
    END
  END Data_Out[4]
  PIN Data_Out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1778.450 0.000 1778.730 4.000 ;
    END
  END Data_Out[5]
  PIN Data_Out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1874.590 0.000 1874.870 4.000 ;
    END
  END Data_Out[6]
  PIN Data_Out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1970.730 0.000 1971.010 4.000 ;
    END
  END Data_Out[7]
  PIN PreCharge
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1249.910 2996.000 1250.190 3000.000 ;
    END
  END PreCharge
  PIN Proj_Select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END Proj_Select[0]
  PIN Proj_Select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1165.560 4.000 1166.160 ;
    END
  END Proj_Select[1]
  PIN ReadEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END ReadEnable
  PIN Reram_In_Enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2831.560 4.000 2832.160 ;
    END
  END Reram_In_Enable
  PIN Trunc_Enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2165.160 4.000 2165.760 ;
    END
  END Trunc_Enable
  PIN WL_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END WL_enable
  PIN WriteEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END WriteEnable
  PIN analog_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.430 0.000 2451.710 4.000 ;
    END
  END analog_io1
  PIN analog_io2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2498.360 4.000 2498.960 ;
    END
  END analog_io2
  PIN analog_io3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.290 0.000 2355.570 4.000 ;
    END
  END analog_io3
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 975.160 2500.000 975.760 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2471.160 2500.000 2471.760 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2620.760 2500.000 2621.360 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2770.360 2500.000 2770.960 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2919.960 2500.000 2920.560 ;
    END
  END io_oeb[13]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1124.760 2500.000 1125.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1274.360 2500.000 1274.960 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1423.960 2500.000 1424.560 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1573.560 2500.000 1574.160 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1723.160 2500.000 1723.760 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1872.760 2500.000 1873.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2022.360 2500.000 2022.960 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2171.960 2500.000 2172.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2321.560 2500.000 2322.160 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 77.560 2500.000 78.160 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 227.160 2500.000 227.760 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 376.760 2500.000 377.360 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 526.360 2500.000 526.960 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 675.960 2500.000 676.560 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 825.560 2500.000 826.160 ;
    END
  END io_out[5]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END rst
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.870 0.000 2067.150 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.010 0.000 2163.290 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2259.150 0.000 2259.430 4.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 958.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 981.800 2019.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 2986.800 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 72.240 10.640 73.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.840 10.640 227.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 379.440 10.640 381.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.040 10.640 534.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 686.640 10.640 688.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 840.240 10.640 841.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 993.840 10.640 995.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.440 10.640 1149.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.040 10.640 1302.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.640 10.640 1456.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.240 10.640 1609.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1761.840 10.640 1763.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1915.440 10.640 1917.040 958.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1915.440 981.800 1917.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2069.040 10.640 2070.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2222.640 10.640 2224.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.240 10.640 2377.840 2986.800 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 123.440 10.640 125.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.040 10.640 278.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 430.640 10.640 432.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.240 10.640 585.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 737.840 10.640 739.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.440 10.640 893.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1045.040 10.640 1046.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.640 10.640 1200.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1352.240 10.640 1353.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1505.840 10.640 1507.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1659.440 10.640 1661.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1813.040 10.640 1814.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.640 10.640 1968.240 958.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.640 981.800 1968.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2120.240 10.640 2121.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2273.840 10.640 2275.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2427.440 10.640 2429.040 2986.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 149.040 10.640 150.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 302.640 10.640 304.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.240 10.640 457.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 609.840 10.640 611.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 763.440 10.640 765.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.040 10.640 918.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1070.640 10.640 1072.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.240 10.640 1225.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.840 10.640 1379.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.440 10.640 1533.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1685.040 10.640 1686.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1838.640 10.640 1840.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1992.240 10.640 1993.840 958.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1992.240 981.800 1993.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.840 10.640 2147.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2299.440 10.640 2301.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2453.040 10.640 2454.640 2986.800 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.640 10.640 48.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.240 10.640 201.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.840 10.640 355.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.440 10.640 509.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.040 10.640 662.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.640 10.640 816.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 968.240 10.640 969.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.840 10.640 1123.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.440 10.640 1277.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1429.040 10.640 1430.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1582.640 10.640 1584.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.240 10.640 1737.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1889.840 10.640 1891.440 958.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1889.840 981.800 1891.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2043.440 10.640 2045.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.040 10.640 2198.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2350.640 10.640 2352.240 2986.800 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 958.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 981.800 1942.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 2986.800 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2494.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 2494.120 2986.800 ;
      LAYER met2 ;
        RECT 4.690 2995.720 1249.630 2996.000 ;
        RECT 1250.470 2995.720 2493.570 2996.000 ;
        RECT 4.690 4.280 2493.570 2995.720 ;
        RECT 4.690 3.670 47.650 4.280 ;
        RECT 48.490 3.670 143.790 4.280 ;
        RECT 144.630 3.670 239.930 4.280 ;
        RECT 240.770 3.670 336.070 4.280 ;
        RECT 336.910 3.670 432.210 4.280 ;
        RECT 433.050 3.670 528.350 4.280 ;
        RECT 529.190 3.670 624.490 4.280 ;
        RECT 625.330 3.670 720.630 4.280 ;
        RECT 721.470 3.670 816.770 4.280 ;
        RECT 817.610 3.670 912.910 4.280 ;
        RECT 913.750 3.670 1009.050 4.280 ;
        RECT 1009.890 3.670 1105.190 4.280 ;
        RECT 1106.030 3.670 1201.330 4.280 ;
        RECT 1202.170 3.670 1297.470 4.280 ;
        RECT 1298.310 3.670 1393.610 4.280 ;
        RECT 1394.450 3.670 1489.750 4.280 ;
        RECT 1490.590 3.670 1585.890 4.280 ;
        RECT 1586.730 3.670 1682.030 4.280 ;
        RECT 1682.870 3.670 1778.170 4.280 ;
        RECT 1779.010 3.670 1874.310 4.280 ;
        RECT 1875.150 3.670 1970.450 4.280 ;
        RECT 1971.290 3.670 2066.590 4.280 ;
        RECT 2067.430 3.670 2162.730 4.280 ;
        RECT 2163.570 3.670 2258.870 4.280 ;
        RECT 2259.710 3.670 2355.010 4.280 ;
        RECT 2355.850 3.670 2451.150 4.280 ;
        RECT 2451.990 3.670 2493.570 4.280 ;
      LAYER met3 ;
        RECT 4.000 2920.960 2496.000 2986.725 ;
        RECT 4.000 2919.560 2495.600 2920.960 ;
        RECT 4.000 2832.560 2496.000 2919.560 ;
        RECT 4.400 2831.160 2496.000 2832.560 ;
        RECT 4.000 2771.360 2496.000 2831.160 ;
        RECT 4.000 2769.960 2495.600 2771.360 ;
        RECT 4.000 2621.760 2496.000 2769.960 ;
        RECT 4.000 2620.360 2495.600 2621.760 ;
        RECT 4.000 2499.360 2496.000 2620.360 ;
        RECT 4.400 2497.960 2496.000 2499.360 ;
        RECT 4.000 2472.160 2496.000 2497.960 ;
        RECT 4.000 2470.760 2495.600 2472.160 ;
        RECT 4.000 2322.560 2496.000 2470.760 ;
        RECT 4.000 2321.160 2495.600 2322.560 ;
        RECT 4.000 2172.960 2496.000 2321.160 ;
        RECT 4.000 2171.560 2495.600 2172.960 ;
        RECT 4.000 2166.160 2496.000 2171.560 ;
        RECT 4.400 2164.760 2496.000 2166.160 ;
        RECT 4.000 2023.360 2496.000 2164.760 ;
        RECT 4.000 2021.960 2495.600 2023.360 ;
        RECT 4.000 1873.760 2496.000 2021.960 ;
        RECT 4.000 1872.360 2495.600 1873.760 ;
        RECT 4.000 1832.960 2496.000 1872.360 ;
        RECT 4.400 1831.560 2496.000 1832.960 ;
        RECT 4.000 1724.160 2496.000 1831.560 ;
        RECT 4.000 1722.760 2495.600 1724.160 ;
        RECT 4.000 1574.560 2496.000 1722.760 ;
        RECT 4.000 1573.160 2495.600 1574.560 ;
        RECT 4.000 1499.760 2496.000 1573.160 ;
        RECT 4.400 1498.360 2496.000 1499.760 ;
        RECT 4.000 1424.960 2496.000 1498.360 ;
        RECT 4.000 1423.560 2495.600 1424.960 ;
        RECT 4.000 1275.360 2496.000 1423.560 ;
        RECT 4.000 1273.960 2495.600 1275.360 ;
        RECT 4.000 1166.560 2496.000 1273.960 ;
        RECT 4.400 1165.160 2496.000 1166.560 ;
        RECT 4.000 1125.760 2496.000 1165.160 ;
        RECT 4.000 1124.360 2495.600 1125.760 ;
        RECT 4.000 976.160 2496.000 1124.360 ;
        RECT 4.000 974.760 2495.600 976.160 ;
        RECT 4.000 833.360 2496.000 974.760 ;
        RECT 4.400 831.960 2496.000 833.360 ;
        RECT 4.000 826.560 2496.000 831.960 ;
        RECT 4.000 825.160 2495.600 826.560 ;
        RECT 4.000 676.960 2496.000 825.160 ;
        RECT 4.000 675.560 2495.600 676.960 ;
        RECT 4.000 527.360 2496.000 675.560 ;
        RECT 4.000 525.960 2495.600 527.360 ;
        RECT 4.000 500.160 2496.000 525.960 ;
        RECT 4.400 498.760 2496.000 500.160 ;
        RECT 4.000 377.760 2496.000 498.760 ;
        RECT 4.000 376.360 2495.600 377.760 ;
        RECT 4.000 228.160 2496.000 376.360 ;
        RECT 4.000 226.760 2495.600 228.160 ;
        RECT 4.000 166.960 2496.000 226.760 ;
        RECT 4.400 165.560 2496.000 166.960 ;
        RECT 4.000 78.560 2496.000 165.560 ;
        RECT 4.000 77.160 2495.600 78.560 ;
        RECT 4.000 10.715 2496.000 77.160 ;
      LAYER met4 ;
        RECT 1585.455 13.095 1607.840 2898.665 ;
        RECT 1610.240 13.095 1633.440 2898.665 ;
        RECT 1635.840 13.095 1659.040 2898.665 ;
        RECT 1661.440 13.095 1684.640 2898.665 ;
        RECT 1687.040 13.095 1710.240 2898.665 ;
        RECT 1712.640 13.095 1735.840 2898.665 ;
        RECT 1738.240 13.095 1761.440 2898.665 ;
        RECT 1763.840 13.095 1787.040 2898.665 ;
        RECT 1789.440 13.095 1812.640 2898.665 ;
        RECT 1815.040 13.095 1838.240 2898.665 ;
        RECT 1840.640 13.095 1863.840 2898.665 ;
        RECT 1866.240 981.400 1889.440 2898.665 ;
        RECT 1891.840 981.400 1915.040 2898.665 ;
        RECT 1917.440 981.400 1940.640 2898.665 ;
        RECT 1943.040 981.400 1966.240 2898.665 ;
        RECT 1968.640 981.400 1991.840 2898.665 ;
        RECT 1994.240 981.400 2017.440 2898.665 ;
        RECT 2019.840 981.400 2024.850 2898.665 ;
        RECT 1866.240 958.400 2024.850 981.400 ;
        RECT 1866.240 13.095 1889.440 958.400 ;
        RECT 1891.840 13.095 1915.040 958.400 ;
        RECT 1917.440 13.095 1940.640 958.400 ;
        RECT 1943.040 13.095 1966.240 958.400 ;
        RECT 1968.640 13.095 1991.840 958.400 ;
        RECT 1994.240 13.095 2017.440 958.400 ;
        RECT 2019.840 13.095 2024.850 958.400 ;
  END
END user_proj_IMPACT_HEAD
END LIBRARY

